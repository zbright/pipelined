`include "register_file_if.vh"
`include "cpu_types_pkg.vh"

module register_file (
	input logic CLK,
	input logic nRST,
	register_file_if.rf registerval
	);
	
	logic [31:0] [31:0] storeregister; 
	logic [2:0] k;	

	always_ff @(negedge CLK, negedge nRST)
		begin: WRITE
			if (nRST == 0) begin
				storeregister <= '0;
			end else if (registerval.WEN) begin
				if (registerval.wsel) begin
					storeregister[registerval.wsel] <= registerval.wdat;
				end else if (registerval.wsel == 0) begin
					storeregister[0] <= 0;
				end
			end
		end

	always_comb
		begin
			registerval.rdat1 = storeregister[registerval.rsel1];
			registerval.rdat2 = storeregister[registerval.rsel2];
		end
		
endmodule	
	


	
	

