// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 32-bit"
// VERSION "Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"

// DATE "03/06/2014 12:16:32"

// 
// Device: Altera EP4CE115F29C8 Package FBGA780
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	CLK,
	nRST,
	\syif.halt ,
	\syif.load ,
	\syif.addr ,
	\syif.store ,
	\syif.REN ,
	\syif.WEN ,
	\syif.tbCTRL );
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	CLK;
input 	nRST;
output 	\syif.halt ;
output 	[31:0] \syif.load ;
input 	[31:0] \syif.addr ;
input 	[31:0] \syif.store ;
input 	\syif.REN ;
input 	\syif.WEN ;
input 	\syif.tbCTRL ;

// Design Ports Information
// syif.halt	=>  Location: PIN_D15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[0]	=>  Location: PIN_D14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[1]	=>  Location: PIN_P1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[2]	=>  Location: PIN_AC15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[3]	=>  Location: PIN_P25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[4]	=>  Location: PIN_AA15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[5]	=>  Location: PIN_AC14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[6]	=>  Location: PIN_E25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[7]	=>  Location: PIN_H21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[8]	=>  Location: PIN_G21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[9]	=>  Location: PIN_AC17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[10]	=>  Location: PIN_M23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[11]	=>  Location: PIN_E17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[12]	=>  Location: PIN_C17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[13]	=>  Location: PIN_A19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[14]	=>  Location: PIN_C16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[15]	=>  Location: PIN_C12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[16]	=>  Location: PIN_D13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[17]	=>  Location: PIN_AD11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[18]	=>  Location: PIN_A12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[19]	=>  Location: PIN_AA12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[20]	=>  Location: PIN_AB14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[21]	=>  Location: PIN_AF14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[22]	=>  Location: PIN_Y13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[23]	=>  Location: PIN_G14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[24]	=>  Location: PIN_AA13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[25]	=>  Location: PIN_C13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[26]	=>  Location: PIN_AG12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[27]	=>  Location: PIN_AH12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[28]	=>  Location: PIN_B19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[29]	=>  Location: PIN_AG17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[30]	=>  Location: PIN_AD15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[31]	=>  Location: PIN_Y15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.WEN	=>  Location: PIN_AG15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.tbCTRL	=>  Location: PIN_AH15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.REN	=>  Location: PIN_AE15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[0]	=>  Location: PIN_D16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[1]	=>  Location: PIN_Y12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[3]	=>  Location: PIN_H15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[2]	=>  Location: PIN_H17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[5]	=>  Location: PIN_D12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[4]	=>  Location: PIN_P2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[7]	=>  Location: PIN_C14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[6]	=>  Location: PIN_E15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[9]	=>  Location: PIN_AA14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[8]	=>  Location: PIN_J15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[11]	=>  Location: PIN_P27,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[10]	=>  Location: PIN_N21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[13]	=>  Location: PIN_AH17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[12]	=>  Location: PIN_G16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[15]	=>  Location: PIN_AD14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[14]	=>  Location: PIN_F15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[17]	=>  Location: PIN_G18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[16]	=>  Location: PIN_H16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[19]	=>  Location: PIN_AF17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[18]	=>  Location: PIN_G19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[21]	=>  Location: PIN_AE17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[20]	=>  Location: PIN_AB15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[23]	=>  Location: PIN_B17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[22]	=>  Location: PIN_J14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[25]	=>  Location: PIN_L1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[24]	=>  Location: PIN_L2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[27]	=>  Location: PIN_Y14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[26]	=>  Location: PIN_H14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[29]	=>  Location: PIN_P28,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[28]	=>  Location: PIN_F14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[31]	=>  Location: PIN_A17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[30]	=>  Location: PIN_C15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// nRST	=>  Location: PIN_Y2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// CLK	=>  Location: PIN_J1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[0]	=>  Location: PIN_AH21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[1]	=>  Location: PIN_J19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[2]	=>  Location: PIN_J16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[3]	=>  Location: PIN_AC11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[4]	=>  Location: PIN_G15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[5]	=>  Location: PIN_AD17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[6]	=>  Location: PIN_J17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[7]	=>  Location: PIN_P21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[8]	=>  Location: PIN_F17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[9]	=>  Location: PIN_R27,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[10]	=>  Location: PIN_R22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[11]	=>  Location: PIN_AG18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[12]	=>  Location: PIN_A18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[13]	=>  Location: PIN_AH19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[14]	=>  Location: PIN_AG19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[15]	=>  Location: PIN_G22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[16]	=>  Location: PIN_R24,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[17]	=>  Location: PIN_R7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[18]	=>  Location: PIN_R21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[19]	=>  Location: PIN_H19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[20]	=>  Location: PIN_AA16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[21]	=>  Location: PIN_R28,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[22]	=>  Location: PIN_AF15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[23]	=>  Location: PIN_AE14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[24]	=>  Location: PIN_AF16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[25]	=>  Location: PIN_G20,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[26]	=>  Location: PIN_AH18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[27]	=>  Location: PIN_R25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[28]	=>  Location: PIN_B18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[29]	=>  Location: PIN_AB16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[30]	=>  Location: PIN_AG21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[31]	=>  Location: PIN_AE16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tms	=>  Location: PIN_P8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tck	=>  Location: PIN_P5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdi	=>  Location: PIN_P7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdo	=>  Location: PIN_P6,	 I/O Standard: 2.5 V,	 Current Strength: Default


wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ;
wire \CPU|DP|dpif.halt~q ;
wire \CPU|DP|EXMEM|temp_dmemWEN~q ;
wire \CPU|DP|EXMEM|temp_dmemREN~q ;
wire \ramaddr~0_combout ;
wire \ramaddr~1_combout ;
wire \ramaddr~2_combout ;
wire \ramaddr~3_combout ;
wire \ramaddr~4_combout ;
wire \ramaddr~5_combout ;
wire \ramaddr~6_combout ;
wire \ramaddr~7_combout ;
wire \ramaddr~8_combout ;
wire \ramaddr~9_combout ;
wire \ramaddr~10_combout ;
wire \ramaddr~11_combout ;
wire \ramaddr~12_combout ;
wire \ramaddr~13_combout ;
wire \ramaddr~14_combout ;
wire \ramaddr~15_combout ;
wire \ramaddr~16_combout ;
wire \ramaddr~17_combout ;
wire \ramaddr~18_combout ;
wire \ramaddr~19_combout ;
wire \ramaddr~20_combout ;
wire \ramaddr~21_combout ;
wire \ramaddr~22_combout ;
wire \ramaddr~23_combout ;
wire \ramaddr~24_combout ;
wire \ramaddr~25_combout ;
wire \ramaddr~26_combout ;
wire \ramaddr~27_combout ;
wire \ramaddr~28_combout ;
wire \ramaddr~29_combout ;
wire \ramaddr~30_combout ;
wire \ramaddr~31_combout ;
wire \ramaddr~32_combout ;
wire \ramaddr~33_combout ;
wire \ramaddr~34_combout ;
wire \ramaddr~35_combout ;
wire \ramaddr~36_combout ;
wire \ramaddr~37_combout ;
wire \ramaddr~38_combout ;
wire \ramaddr~39_combout ;
wire \ramaddr~40_combout ;
wire \ramaddr~41_combout ;
wire \ramaddr~42_combout ;
wire \ramaddr~43_combout ;
wire \ramaddr~44_combout ;
wire \ramaddr~45_combout ;
wire \ramaddr~46_combout ;
wire \ramaddr~47_combout ;
wire \ramaddr~48_combout ;
wire \ramaddr~49_combout ;
wire \ramaddr~50_combout ;
wire \ramaddr~51_combout ;
wire \ramaddr~52_combout ;
wire \ramaddr~53_combout ;
wire \ramaddr~54_combout ;
wire \ramaddr~55_combout ;
wire \RAM|always1~2_combout ;
wire \RAM|ramif.ramload[0]~0_combout ;
wire \RAM|ramif.ramload[1]~1_combout ;
wire \RAM|ramif.ramload[2]~2_combout ;
wire \RAM|ramif.ramload[3]~3_combout ;
wire \RAM|ramif.ramload[4]~4_combout ;
wire \RAM|ramif.ramload[5]~5_combout ;
wire \RAM|ramif.ramload[6]~6_combout ;
wire \RAM|ramif.ramload[7]~7_combout ;
wire \RAM|ramif.ramload[8]~8_combout ;
wire \RAM|ramif.ramload[9]~9_combout ;
wire \RAM|ramif.ramload[10]~10_combout ;
wire \RAM|ramif.ramload[11]~11_combout ;
wire \RAM|ramif.ramload[12]~12_combout ;
wire \RAM|ramif.ramload[13]~13_combout ;
wire \RAM|ramif.ramload[14]~14_combout ;
wire \RAM|ramif.ramload[15]~15_combout ;
wire \RAM|ramif.ramload[16]~16_combout ;
wire \RAM|ramif.ramload[17]~17_combout ;
wire \RAM|ramif.ramload[18]~18_combout ;
wire \RAM|ramif.ramload[19]~19_combout ;
wire \RAM|ramif.ramload[20]~20_combout ;
wire \RAM|ramif.ramload[21]~21_combout ;
wire \RAM|ramif.ramload[22]~22_combout ;
wire \RAM|ramif.ramload[23]~23_combout ;
wire \RAM|ramif.ramload[24]~24_combout ;
wire \RAM|ramif.ramload[25]~25_combout ;
wire \RAM|ramif.ramload[26]~26_combout ;
wire \RAM|ramif.ramload[27]~27_combout ;
wire \RAM|ramif.ramload[28]~28_combout ;
wire \RAM|ramif.ramload[29]~29_combout ;
wire \RAM|ramif.ramload[30]~30_combout ;
wire \RAM|ramif.ramload[31]~31_combout ;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ;
wire \CPUCLK~q ;
wire \ramWEN~0_combout ;
wire \ramWEN~1_combout ;
wire \ramstore~0_combout ;
wire \ramaddr~56_combout ;
wire \ramaddr~57_combout ;
wire \ramaddr~58_combout ;
wire \ramaddr~59_combout ;
wire \ramaddr~60_combout ;
wire \ramaddr~61_combout ;
wire \ramaddr~62_combout ;
wire \ramaddr~63_combout ;
wire \ramstore~1_combout ;
wire \ramstore~2_combout ;
wire \ramstore~3_combout ;
wire \ramstore~4_combout ;
wire \ramstore~5_combout ;
wire \ramstore~6_combout ;
wire \ramstore~7_combout ;
wire \ramstore~8_combout ;
wire \ramstore~9_combout ;
wire \ramstore~10_combout ;
wire \ramstore~11_combout ;
wire \ramstore~12_combout ;
wire \ramstore~13_combout ;
wire \ramstore~14_combout ;
wire \ramstore~15_combout ;
wire \ramstore~16_combout ;
wire \ramstore~17_combout ;
wire \ramstore~18_combout ;
wire \ramstore~19_combout ;
wire \ramstore~20_combout ;
wire \ramstore~21_combout ;
wire \ramstore~22_combout ;
wire \ramstore~23_combout ;
wire \ramstore~24_combout ;
wire \ramstore~25_combout ;
wire \ramstore~26_combout ;
wire \ramstore~27_combout ;
wire \ramstore~28_combout ;
wire \ramstore~29_combout ;
wire \ramstore~30_combout ;
wire \ramstore~31_combout ;
wire \Equal0~0_combout ;
wire \CPUCLK~0_combout ;
wire \ramREN~0_combout ;
wire \count[3]~0_combout ;
wire \count[2]~1_combout ;
wire \count[1]~2_combout ;
wire \count~3_combout ;
wire \ramaddr~25_wirecell_combout ;
wire \altera_internal_jtag~TCKUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ;
wire \syif.WEN~input_o ;
wire \syif.tbCTRL~input_o ;
wire \syif.REN~input_o ;
wire \syif.addr[0]~input_o ;
wire \syif.addr[1]~input_o ;
wire \syif.addr[3]~input_o ;
wire \syif.addr[2]~input_o ;
wire \syif.addr[5]~input_o ;
wire \syif.addr[4]~input_o ;
wire \syif.addr[7]~input_o ;
wire \syif.addr[6]~input_o ;
wire \syif.addr[9]~input_o ;
wire \syif.addr[8]~input_o ;
wire \syif.addr[11]~input_o ;
wire \syif.addr[10]~input_o ;
wire \syif.addr[13]~input_o ;
wire \syif.addr[12]~input_o ;
wire \syif.addr[15]~input_o ;
wire \syif.addr[14]~input_o ;
wire \syif.addr[17]~input_o ;
wire \syif.addr[16]~input_o ;
wire \syif.addr[19]~input_o ;
wire \syif.addr[18]~input_o ;
wire \syif.addr[21]~input_o ;
wire \syif.addr[20]~input_o ;
wire \syif.addr[23]~input_o ;
wire \syif.addr[22]~input_o ;
wire \syif.addr[25]~input_o ;
wire \syif.addr[24]~input_o ;
wire \syif.addr[27]~input_o ;
wire \syif.addr[26]~input_o ;
wire \syif.addr[29]~input_o ;
wire \syif.addr[28]~input_o ;
wire \syif.addr[31]~input_o ;
wire \syif.addr[30]~input_o ;
wire \nRST~input_o ;
wire \CLK~input_o ;
wire \syif.store[0]~input_o ;
wire \syif.store[1]~input_o ;
wire \syif.store[2]~input_o ;
wire \syif.store[3]~input_o ;
wire \syif.store[4]~input_o ;
wire \syif.store[5]~input_o ;
wire \syif.store[6]~input_o ;
wire \syif.store[7]~input_o ;
wire \syif.store[8]~input_o ;
wire \syif.store[9]~input_o ;
wire \syif.store[10]~input_o ;
wire \syif.store[11]~input_o ;
wire \syif.store[12]~input_o ;
wire \syif.store[13]~input_o ;
wire \syif.store[14]~input_o ;
wire \syif.store[15]~input_o ;
wire \syif.store[16]~input_o ;
wire \syif.store[17]~input_o ;
wire \syif.store[18]~input_o ;
wire \syif.store[19]~input_o ;
wire \syif.store[20]~input_o ;
wire \syif.store[21]~input_o ;
wire \syif.store[22]~input_o ;
wire \syif.store[23]~input_o ;
wire \syif.store[24]~input_o ;
wire \syif.store[25]~input_o ;
wire \syif.store[26]~input_o ;
wire \syif.store[27]~input_o ;
wire \syif.store[28]~input_o ;
wire \syif.store[29]~input_o ;
wire \syif.store[30]~input_o ;
wire \syif.store[31]~input_o ;
wire \altera_internal_jtag~TCKUTAPclkctrl_outclk ;
wire \CPUCLK~clkctrl_outclk ;
wire \nRST~inputclkctrl_outclk ;
wire \CLK~inputclkctrl_outclk ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ;
wire \~QIC_CREATED_GND~I_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg ;
wire [9:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg ;
wire [5:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt ;
wire [15:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR ;
wire [3:0] count;
wire [31:0] \CPU|DP|PC|pccount ;
wire [3:0] \RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg ;
wire [31:0] \CPU|DP|EXMEM|temp_rdat2 ;
wire [31:0] \CPU|DP|EXMEM|temp_aluResult ;


ram RAM(
	.is_in_use_reg(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.temp_dmemWEN(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.temp_dmemREN(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.ramaddr(\ramaddr~0_combout ),
	.ramaddr1(\ramaddr~1_combout ),
	.ramaddr2(\ramaddr~2_combout ),
	.ramaddr3(\ramaddr~3_combout ),
	.ramaddr4(\ramaddr~5_combout ),
	.ramaddr5(\ramaddr~7_combout ),
	.ramaddr6(\ramaddr~9_combout ),
	.ramaddr7(\ramaddr~11_combout ),
	.ramaddr8(\ramaddr~13_combout ),
	.ramaddr9(\ramaddr~15_combout ),
	.ramaddr10(\ramaddr~17_combout ),
	.ramaddr11(\ramaddr~19_combout ),
	.ramaddr12(\ramaddr~21_combout ),
	.ramaddr13(\ramaddr~23_combout ),
	.ramaddr14(\ramaddr~25_combout ),
	.ramaddr15(\ramaddr~27_combout ),
	.\ramif.ramaddr ({\ramaddr~53_combout ,\ramaddr~55_combout ,\ramaddr~49_combout ,\ramaddr~51_combout ,\ramaddr~62_combout ,\ramaddr~63_combout ,\ramaddr~43_combout ,\ramaddr~45_combout ,\ramaddr~39_combout ,gnd,\ramaddr~60_combout ,\ramaddr~61_combout ,\ramaddr~33_combout ,
\ramaddr~35_combout ,\ramaddr~29_combout ,\ramaddr~31_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\ramaddr~59_combout ,\ramaddr~58_combout }),
	.ramaddr16(\ramaddr~36_combout ),
	.ramaddr17(\ramaddr~37_combout ),
	.ramaddr18(\ramaddr~41_combout ),
	.ramaddr19(\ramaddr~46_combout ),
	.ramaddr20(\ramaddr~47_combout ),
	.always1(\RAM|always1~2_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~16_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~17_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~18_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~19_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~20_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~21_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~22_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~23_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~24_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~25_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~26_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~27_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~28_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~29_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~30_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~31_combout ),
	.ir_loaded_address_reg_0(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.ir_loaded_address_reg_1(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.ir_loaded_address_reg_2(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.ir_loaded_address_reg_3(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.tdo(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.ramWEN(\ramWEN~0_combout ),
	.ramstore(\ramstore~0_combout ),
	.ramaddr21(\ramaddr~56_combout ),
	.ramaddr22(\ramaddr~57_combout ),
	.ramstore1(\ramstore~1_combout ),
	.ramstore2(\ramstore~2_combout ),
	.ramstore3(\ramstore~3_combout ),
	.ramstore4(\ramstore~4_combout ),
	.ramstore5(\ramstore~5_combout ),
	.ramstore6(\ramstore~6_combout ),
	.ramstore7(\ramstore~7_combout ),
	.ramstore8(\ramstore~8_combout ),
	.ramstore9(\ramstore~9_combout ),
	.ramstore10(\ramstore~10_combout ),
	.ramstore11(\ramstore~11_combout ),
	.ramstore12(\ramstore~12_combout ),
	.ramstore13(\ramstore~13_combout ),
	.ramstore14(\ramstore~14_combout ),
	.ramstore15(\ramstore~15_combout ),
	.ramstore16(\ramstore~16_combout ),
	.ramstore17(\ramstore~17_combout ),
	.ramstore18(\ramstore~18_combout ),
	.ramstore19(\ramstore~19_combout ),
	.ramstore20(\ramstore~20_combout ),
	.ramstore21(\ramstore~21_combout ),
	.ramstore22(\ramstore~22_combout ),
	.ramstore23(\ramstore~23_combout ),
	.ramstore24(\ramstore~24_combout ),
	.ramstore25(\ramstore~25_combout ),
	.ramstore26(\ramstore~26_combout ),
	.ramstore27(\ramstore~27_combout ),
	.ramstore28(\ramstore~28_combout ),
	.ramstore29(\ramstore~29_combout ),
	.ramstore30(\ramstore~30_combout ),
	.ramstore31(\ramstore~31_combout ),
	.\ramif.ramREN (\ramREN~0_combout ),
	.ramaddr23(\ramaddr~25_wirecell_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.irf_reg_0_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.irf_reg_2_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.irf_reg_3_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.irf_reg_4_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.node_ena_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.clr_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.virtual_ir_scan_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.state_5(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.state_8(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.syifWEN(\syif.WEN~input_o ),
	.syiftbCTRL(\syif.tbCTRL~input_o ),
	.syifREN(\syif.REN~input_o ),
	.syifaddr_0(\syif.addr[0]~input_o ),
	.syifaddr_1(\syif.addr[1]~input_o ),
	.syifaddr_3(\syif.addr[3]~input_o ),
	.syifaddr_2(\syif.addr[2]~input_o ),
	.syifaddr_21(\syif.addr[21]~input_o ),
	.syifaddr_20(\syif.addr[20]~input_o ),
	.syifaddr_27(\syif.addr[27]~input_o ),
	.syifaddr_26(\syif.addr[26]~input_o ),
	.nRST(\nRST~input_o ),
	.altera_internal_jtag1(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.CLK(\CLK~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pipeline CPU(
	.dpifhalt(\CPU|DP|dpif.halt~q ),
	.temp_aluResult_1(\CPU|DP|EXMEM|temp_aluResult [1]),
	.pccount_1(\CPU|DP|PC|pccount [1]),
	.temp_dmemWEN(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.temp_dmemREN(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.temp_aluResult_0(\CPU|DP|EXMEM|temp_aluResult [0]),
	.pccount_0(\CPU|DP|PC|pccount [0]),
	.temp_aluResult_2(\CPU|DP|EXMEM|temp_aluResult [2]),
	.pccount_2(\CPU|DP|PC|pccount [2]),
	.temp_aluResult_3(\CPU|DP|EXMEM|temp_aluResult [3]),
	.pccount_3(\CPU|DP|PC|pccount [3]),
	.temp_aluResult_5(\CPU|DP|EXMEM|temp_aluResult [5]),
	.pccount_5(\CPU|DP|PC|pccount [5]),
	.temp_aluResult_4(\CPU|DP|EXMEM|temp_aluResult [4]),
	.pccount_4(\CPU|DP|PC|pccount [4]),
	.temp_aluResult_7(\CPU|DP|EXMEM|temp_aluResult [7]),
	.pccount_7(\CPU|DP|PC|pccount [7]),
	.temp_aluResult_6(\CPU|DP|EXMEM|temp_aluResult [6]),
	.pccount_6(\CPU|DP|PC|pccount [6]),
	.temp_aluResult_9(\CPU|DP|EXMEM|temp_aluResult [9]),
	.pccount_9(\CPU|DP|PC|pccount [9]),
	.temp_aluResult_8(\CPU|DP|EXMEM|temp_aluResult [8]),
	.pccount_8(\CPU|DP|PC|pccount [8]),
	.temp_aluResult_11(\CPU|DP|EXMEM|temp_aluResult [11]),
	.pccount_11(\CPU|DP|PC|pccount [11]),
	.temp_aluResult_10(\CPU|DP|EXMEM|temp_aluResult [10]),
	.pccount_10(\CPU|DP|PC|pccount [10]),
	.temp_aluResult_13(\CPU|DP|EXMEM|temp_aluResult [13]),
	.pccount_13(\CPU|DP|PC|pccount [13]),
	.temp_aluResult_12(\CPU|DP|EXMEM|temp_aluResult [12]),
	.pccount_12(\CPU|DP|PC|pccount [12]),
	.temp_aluResult_15(\CPU|DP|EXMEM|temp_aluResult [15]),
	.pccount_15(\CPU|DP|PC|pccount [15]),
	.temp_aluResult_14(\CPU|DP|EXMEM|temp_aluResult [14]),
	.pccount_14(\CPU|DP|PC|pccount [14]),
	.temp_aluResult_17(\CPU|DP|EXMEM|temp_aluResult [17]),
	.pccount_17(\CPU|DP|PC|pccount [17]),
	.temp_aluResult_16(\CPU|DP|EXMEM|temp_aluResult [16]),
	.pccount_16(\CPU|DP|PC|pccount [16]),
	.temp_aluResult_19(\CPU|DP|EXMEM|temp_aluResult [19]),
	.pccount_19(\CPU|DP|PC|pccount [19]),
	.temp_aluResult_18(\CPU|DP|EXMEM|temp_aluResult [18]),
	.pccount_18(\CPU|DP|PC|pccount [18]),
	.temp_aluResult_20(\CPU|DP|EXMEM|temp_aluResult [20]),
	.pccount_20(\CPU|DP|PC|pccount [20]),
	.temp_aluResult_21(\CPU|DP|EXMEM|temp_aluResult [21]),
	.pccount_21(\CPU|DP|PC|pccount [21]),
	.temp_aluResult_23(\CPU|DP|EXMEM|temp_aluResult [23]),
	.pccount_23(\CPU|DP|PC|pccount [23]),
	.temp_aluResult_22(\CPU|DP|EXMEM|temp_aluResult [22]),
	.pccount_22(\CPU|DP|PC|pccount [22]),
	.temp_aluResult_25(\CPU|DP|EXMEM|temp_aluResult [25]),
	.pccount_25(\CPU|DP|PC|pccount [25]),
	.temp_aluResult_24(\CPU|DP|EXMEM|temp_aluResult [24]),
	.pccount_24(\CPU|DP|PC|pccount [24]),
	.temp_aluResult_26(\CPU|DP|EXMEM|temp_aluResult [26]),
	.pccount_26(\CPU|DP|PC|pccount [26]),
	.temp_aluResult_27(\CPU|DP|EXMEM|temp_aluResult [27]),
	.pccount_27(\CPU|DP|PC|pccount [27]),
	.temp_aluResult_29(\CPU|DP|EXMEM|temp_aluResult [29]),
	.pccount_29(\CPU|DP|PC|pccount [29]),
	.temp_aluResult_28(\CPU|DP|EXMEM|temp_aluResult [28]),
	.pccount_28(\CPU|DP|PC|pccount [28]),
	.temp_aluResult_31(\CPU|DP|EXMEM|temp_aluResult [31]),
	.pccount_31(\CPU|DP|PC|pccount [31]),
	.temp_aluResult_30(\CPU|DP|EXMEM|temp_aluResult [30]),
	.pccount_30(\CPU|DP|PC|pccount [30]),
	.always1(\RAM|always1~2_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~16_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~17_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~18_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~19_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~20_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~21_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~22_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~23_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~24_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~25_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~26_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~27_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~28_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~29_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~30_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~31_combout ),
	.temp_rdat2_0(\CPU|DP|EXMEM|temp_rdat2 [0]),
	.temp_rdat2_1(\CPU|DP|EXMEM|temp_rdat2 [1]),
	.temp_rdat2_2(\CPU|DP|EXMEM|temp_rdat2 [2]),
	.temp_rdat2_3(\CPU|DP|EXMEM|temp_rdat2 [3]),
	.temp_rdat2_4(\CPU|DP|EXMEM|temp_rdat2 [4]),
	.temp_rdat2_5(\CPU|DP|EXMEM|temp_rdat2 [5]),
	.temp_rdat2_6(\CPU|DP|EXMEM|temp_rdat2 [6]),
	.temp_rdat2_7(\CPU|DP|EXMEM|temp_rdat2 [7]),
	.temp_rdat2_8(\CPU|DP|EXMEM|temp_rdat2 [8]),
	.temp_rdat2_9(\CPU|DP|EXMEM|temp_rdat2 [9]),
	.temp_rdat2_10(\CPU|DP|EXMEM|temp_rdat2 [10]),
	.temp_rdat2_11(\CPU|DP|EXMEM|temp_rdat2 [11]),
	.temp_rdat2_12(\CPU|DP|EXMEM|temp_rdat2 [12]),
	.temp_rdat2_13(\CPU|DP|EXMEM|temp_rdat2 [13]),
	.temp_rdat2_14(\CPU|DP|EXMEM|temp_rdat2 [14]),
	.temp_rdat2_15(\CPU|DP|EXMEM|temp_rdat2 [15]),
	.temp_rdat2_16(\CPU|DP|EXMEM|temp_rdat2 [16]),
	.temp_rdat2_17(\CPU|DP|EXMEM|temp_rdat2 [17]),
	.temp_rdat2_18(\CPU|DP|EXMEM|temp_rdat2 [18]),
	.temp_rdat2_19(\CPU|DP|EXMEM|temp_rdat2 [19]),
	.temp_rdat2_20(\CPU|DP|EXMEM|temp_rdat2 [20]),
	.temp_rdat2_21(\CPU|DP|EXMEM|temp_rdat2 [21]),
	.temp_rdat2_22(\CPU|DP|EXMEM|temp_rdat2 [22]),
	.temp_rdat2_23(\CPU|DP|EXMEM|temp_rdat2 [23]),
	.temp_rdat2_24(\CPU|DP|EXMEM|temp_rdat2 [24]),
	.temp_rdat2_25(\CPU|DP|EXMEM|temp_rdat2 [25]),
	.temp_rdat2_26(\CPU|DP|EXMEM|temp_rdat2 [26]),
	.temp_rdat2_27(\CPU|DP|EXMEM|temp_rdat2 [27]),
	.temp_rdat2_28(\CPU|DP|EXMEM|temp_rdat2 [28]),
	.temp_rdat2_29(\CPU|DP|EXMEM|temp_rdat2 [29]),
	.temp_rdat2_30(\CPU|DP|EXMEM|temp_rdat2 [30]),
	.temp_rdat2_31(\CPU|DP|EXMEM|temp_rdat2 [31]),
	.CPUCLK(\CPUCLK~clkctrl_outclk ),
	.nRST(\nRST~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X63_Y43_N12
cycloneive_lcell_comb \ramaddr~0 (
// Equation(s):
// \ramaddr~0_combout  = (temp_dmemREN1 & (temp_aluResult_1)) # (!temp_dmemREN1 & ((temp_dmemWEN1 & (temp_aluResult_1)) # (!temp_dmemWEN1 & ((pccount_1)))))

	.dataa(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datab(\CPU|DP|EXMEM|temp_aluResult [1]),
	.datac(\CPU|DP|PC|pccount [1]),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~0 .lut_mask = 16'hCCD8;
defparam \ramaddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N28
cycloneive_lcell_comb \ramaddr~1 (
// Equation(s):
// \ramaddr~1_combout  = (temp_dmemWEN1 & (temp_aluResult_0)) # (!temp_dmemWEN1 & ((temp_dmemREN1 & (temp_aluResult_0)) # (!temp_dmemREN1 & ((pccount_0)))))

	.dataa(\CPU|DP|EXMEM|temp_aluResult [0]),
	.datab(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datac(\CPU|DP|PC|pccount [0]),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~1 .lut_mask = 16'hAAB8;
defparam \ramaddr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N20
cycloneive_lcell_comb \ramaddr~2 (
// Equation(s):
// \ramaddr~2_combout  = (temp_dmemREN1 & (((temp_aluResult_2)))) # (!temp_dmemREN1 & ((temp_dmemWEN1 & ((temp_aluResult_2))) # (!temp_dmemWEN1 & (pccount_2))))

	.dataa(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datab(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datac(\CPU|DP|PC|pccount [2]),
	.datad(\CPU|DP|EXMEM|temp_aluResult [2]),
	.cin(gnd),
	.combout(\ramaddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~2 .lut_mask = 16'hFE10;
defparam \ramaddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N12
cycloneive_lcell_comb \ramaddr~3 (
// Equation(s):
// \ramaddr~3_combout  = (temp_dmemWEN1 & (((temp_aluResult_3)))) # (!temp_dmemWEN1 & ((temp_dmemREN1 & ((temp_aluResult_3))) # (!temp_dmemREN1 & (pccount_3))))

	.dataa(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datab(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datac(\CPU|DP|PC|pccount [3]),
	.datad(\CPU|DP|EXMEM|temp_aluResult [3]),
	.cin(gnd),
	.combout(\ramaddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~3 .lut_mask = 16'hFE10;
defparam \ramaddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N28
cycloneive_lcell_comb \ramaddr~4 (
// Equation(s):
// \ramaddr~4_combout  = (temp_dmemREN1 & (((temp_aluResult_5)))) # (!temp_dmemREN1 & ((temp_dmemWEN1 & ((temp_aluResult_5))) # (!temp_dmemWEN1 & (pccount_5))))

	.dataa(\CPU|DP|PC|pccount [5]),
	.datab(\CPU|DP|EXMEM|temp_aluResult [5]),
	.datac(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~4 .lut_mask = 16'hCCCA;
defparam \ramaddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N18
cycloneive_lcell_comb \ramaddr~5 (
// Equation(s):
// \ramaddr~5_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~4_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[5]~input_o ),
	.datad(\ramaddr~4_combout ),
	.cin(gnd),
	.combout(\ramaddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~5 .lut_mask = 16'hF3C0;
defparam \ramaddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N8
cycloneive_lcell_comb \ramaddr~6 (
// Equation(s):
// \ramaddr~6_combout  = (temp_dmemREN1 & (temp_aluResult_4)) # (!temp_dmemREN1 & ((temp_dmemWEN1 & (temp_aluResult_4)) # (!temp_dmemWEN1 & ((pccount_4)))))

	.dataa(\CPU|DP|EXMEM|temp_aluResult [4]),
	.datab(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datac(\CPU|DP|PC|pccount [4]),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~6 .lut_mask = 16'hAAB8;
defparam \ramaddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N4
cycloneive_lcell_comb \ramaddr~7 (
// Equation(s):
// \ramaddr~7_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[4]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~6_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[4]~input_o ),
	.datad(\ramaddr~6_combout ),
	.cin(gnd),
	.combout(\ramaddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~7 .lut_mask = 16'hF3C0;
defparam \ramaddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N18
cycloneive_lcell_comb \ramaddr~8 (
// Equation(s):
// \ramaddr~8_combout  = (temp_dmemREN1 & (temp_aluResult_7)) # (!temp_dmemREN1 & ((temp_dmemWEN1 & (temp_aluResult_7)) # (!temp_dmemWEN1 & ((pccount_7)))))

	.dataa(\CPU|DP|EXMEM|temp_aluResult [7]),
	.datab(\CPU|DP|PC|pccount [7]),
	.datac(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~8 .lut_mask = 16'hAAAC;
defparam \ramaddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N14
cycloneive_lcell_comb \ramaddr~9 (
// Equation(s):
// \ramaddr~9_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[7]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~8_combout )))

	.dataa(\syif.addr[7]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~8_combout ),
	.cin(gnd),
	.combout(\ramaddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~9 .lut_mask = 16'hAFA0;
defparam \ramaddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N10
cycloneive_lcell_comb \ramaddr~10 (
// Equation(s):
// \ramaddr~10_combout  = (temp_dmemREN1 & (temp_aluResult_6)) # (!temp_dmemREN1 & ((temp_dmemWEN1 & (temp_aluResult_6)) # (!temp_dmemWEN1 & ((pccount_6)))))

	.dataa(\CPU|DP|EXMEM|temp_aluResult [6]),
	.datab(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datac(\CPU|DP|PC|pccount [6]),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~10 .lut_mask = 16'hAAB8;
defparam \ramaddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N12
cycloneive_lcell_comb \ramaddr~11 (
// Equation(s):
// \ramaddr~11_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[6]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~10_combout )))

	.dataa(gnd),
	.datab(\syif.addr[6]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~10_combout ),
	.cin(gnd),
	.combout(\ramaddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~11 .lut_mask = 16'hCFC0;
defparam \ramaddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N10
cycloneive_lcell_comb \ramaddr~12 (
// Equation(s):
// \ramaddr~12_combout  = (temp_dmemWEN1 & (((temp_aluResult_9)))) # (!temp_dmemWEN1 & ((temp_dmemREN1 & ((temp_aluResult_9))) # (!temp_dmemREN1 & (pccount_9))))

	.dataa(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datab(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datac(\CPU|DP|PC|pccount [9]),
	.datad(\CPU|DP|EXMEM|temp_aluResult [9]),
	.cin(gnd),
	.combout(\ramaddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~12 .lut_mask = 16'hFE10;
defparam \ramaddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N16
cycloneive_lcell_comb \ramaddr~13 (
// Equation(s):
// \ramaddr~13_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[9]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~12_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[9]~input_o ),
	.datad(\ramaddr~12_combout ),
	.cin(gnd),
	.combout(\ramaddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~13 .lut_mask = 16'hF5A0;
defparam \ramaddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N0
cycloneive_lcell_comb \ramaddr~14 (
// Equation(s):
// \ramaddr~14_combout  = (temp_dmemWEN1 & (((temp_aluResult_8)))) # (!temp_dmemWEN1 & ((temp_dmemREN1 & ((temp_aluResult_8))) # (!temp_dmemREN1 & (pccount_8))))

	.dataa(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datab(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datac(\CPU|DP|PC|pccount [8]),
	.datad(\CPU|DP|EXMEM|temp_aluResult [8]),
	.cin(gnd),
	.combout(\ramaddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~14 .lut_mask = 16'hFE10;
defparam \ramaddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N26
cycloneive_lcell_comb \ramaddr~15 (
// Equation(s):
// \ramaddr~15_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[8]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~14_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[8]~input_o ),
	.datad(\ramaddr~14_combout ),
	.cin(gnd),
	.combout(\ramaddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~15 .lut_mask = 16'hF5A0;
defparam \ramaddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N0
cycloneive_lcell_comb \ramaddr~16 (
// Equation(s):
// \ramaddr~16_combout  = (temp_dmemREN1 & (temp_aluResult_11)) # (!temp_dmemREN1 & ((temp_dmemWEN1 & (temp_aluResult_11)) # (!temp_dmemWEN1 & ((pccount_11)))))

	.dataa(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datab(\CPU|DP|EXMEM|temp_aluResult [11]),
	.datac(\CPU|DP|PC|pccount [11]),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~16 .lut_mask = 16'hCCD8;
defparam \ramaddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N14
cycloneive_lcell_comb \ramaddr~17 (
// Equation(s):
// \ramaddr~17_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~16_combout )))

	.dataa(gnd),
	.datab(\syif.addr[11]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~16_combout ),
	.cin(gnd),
	.combout(\ramaddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~17 .lut_mask = 16'hCFC0;
defparam \ramaddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N6
cycloneive_lcell_comb \ramaddr~18 (
// Equation(s):
// \ramaddr~18_combout  = (temp_dmemREN1 & (temp_aluResult_10)) # (!temp_dmemREN1 & ((temp_dmemWEN1 & (temp_aluResult_10)) # (!temp_dmemWEN1 & ((pccount_10)))))

	.dataa(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datab(\CPU|DP|EXMEM|temp_aluResult [10]),
	.datac(\CPU|DP|PC|pccount [10]),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~18 .lut_mask = 16'hCCD8;
defparam \ramaddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N24
cycloneive_lcell_comb \ramaddr~19 (
// Equation(s):
// \ramaddr~19_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[10]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~18_combout )))

	.dataa(gnd),
	.datab(\syif.addr[10]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~18_combout ),
	.cin(gnd),
	.combout(\ramaddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~19 .lut_mask = 16'hCFC0;
defparam \ramaddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N20
cycloneive_lcell_comb \ramaddr~20 (
// Equation(s):
// \ramaddr~20_combout  = (temp_dmemREN1 & (((temp_aluResult_13)))) # (!temp_dmemREN1 & ((temp_dmemWEN1 & ((temp_aluResult_13))) # (!temp_dmemWEN1 & (pccount_13))))

	.dataa(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datab(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datac(\CPU|DP|PC|pccount [13]),
	.datad(\CPU|DP|EXMEM|temp_aluResult [13]),
	.cin(gnd),
	.combout(\ramaddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~20 .lut_mask = 16'hFE10;
defparam \ramaddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N8
cycloneive_lcell_comb \ramaddr~21 (
// Equation(s):
// \ramaddr~21_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[13]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~20_combout )))

	.dataa(\syif.addr[13]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~20_combout ),
	.cin(gnd),
	.combout(\ramaddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~21 .lut_mask = 16'hAFA0;
defparam \ramaddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N2
cycloneive_lcell_comb \ramaddr~22 (
// Equation(s):
// \ramaddr~22_combout  = (temp_dmemREN1 & (((temp_aluResult_12)))) # (!temp_dmemREN1 & ((temp_dmemWEN1 & ((temp_aluResult_12))) # (!temp_dmemWEN1 & (pccount_12))))

	.dataa(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datab(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datac(\CPU|DP|PC|pccount [12]),
	.datad(\CPU|DP|EXMEM|temp_aluResult [12]),
	.cin(gnd),
	.combout(\ramaddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~22 .lut_mask = 16'hFE10;
defparam \ramaddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N22
cycloneive_lcell_comb \ramaddr~23 (
// Equation(s):
// \ramaddr~23_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[12]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~22_combout )))

	.dataa(\syif.addr[12]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~22_combout ),
	.cin(gnd),
	.combout(\ramaddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~23 .lut_mask = 16'hAFA0;
defparam \ramaddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N2
cycloneive_lcell_comb \ramaddr~24 (
// Equation(s):
// \ramaddr~24_combout  = (temp_dmemREN1 & (((temp_aluResult_15)))) # (!temp_dmemREN1 & ((temp_dmemWEN1 & ((temp_aluResult_15))) # (!temp_dmemWEN1 & (pccount_15))))

	.dataa(\CPU|DP|PC|pccount [15]),
	.datab(\CPU|DP|EXMEM|temp_aluResult [15]),
	.datac(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~24 .lut_mask = 16'hCCCA;
defparam \ramaddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N20
cycloneive_lcell_comb \ramaddr~25 (
// Equation(s):
// \ramaddr~25_combout  = (\syif.tbCTRL~input_o  & (!\syif.addr[15]~input_o )) # (!\syif.tbCTRL~input_o  & ((!\ramaddr~24_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[15]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~24_combout ),
	.cin(gnd),
	.combout(\ramaddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~25 .lut_mask = 16'h2277;
defparam \ramaddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N16
cycloneive_lcell_comb \ramaddr~26 (
// Equation(s):
// \ramaddr~26_combout  = (temp_dmemREN1 & (((temp_aluResult_14)))) # (!temp_dmemREN1 & ((temp_dmemWEN1 & ((temp_aluResult_14))) # (!temp_dmemWEN1 & (pccount_14))))

	.dataa(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datab(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datac(\CPU|DP|PC|pccount [14]),
	.datad(\CPU|DP|EXMEM|temp_aluResult [14]),
	.cin(gnd),
	.combout(\ramaddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~26 .lut_mask = 16'hFE10;
defparam \ramaddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N22
cycloneive_lcell_comb \ramaddr~27 (
// Equation(s):
// \ramaddr~27_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~26_combout )))

	.dataa(gnd),
	.datab(\syif.addr[14]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~26_combout ),
	.cin(gnd),
	.combout(\ramaddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~27 .lut_mask = 16'hCFC0;
defparam \ramaddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N16
cycloneive_lcell_comb \ramaddr~28 (
// Equation(s):
// \ramaddr~28_combout  = (temp_dmemREN1 & (((temp_aluResult_17)))) # (!temp_dmemREN1 & ((temp_dmemWEN1 & ((temp_aluResult_17))) # (!temp_dmemWEN1 & (pccount_17))))

	.dataa(\CPU|DP|PC|pccount [17]),
	.datab(\CPU|DP|EXMEM|temp_aluResult [17]),
	.datac(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~28 .lut_mask = 16'hCCCA;
defparam \ramaddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N8
cycloneive_lcell_comb \ramaddr~29 (
// Equation(s):
// \ramaddr~29_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[17]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~28_combout )))

	.dataa(\syif.addr[17]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~28_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29 .lut_mask = 16'hAFA0;
defparam \ramaddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N18
cycloneive_lcell_comb \ramaddr~30 (
// Equation(s):
// \ramaddr~30_combout  = (temp_dmemREN1 & (temp_aluResult_16)) # (!temp_dmemREN1 & ((temp_dmemWEN1 & (temp_aluResult_16)) # (!temp_dmemWEN1 & ((pccount_16)))))

	.dataa(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datab(\CPU|DP|EXMEM|temp_aluResult [16]),
	.datac(\CPU|DP|PC|pccount [16]),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~30 .lut_mask = 16'hCCD8;
defparam \ramaddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N10
cycloneive_lcell_comb \ramaddr~31 (
// Equation(s):
// \ramaddr~31_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[16]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~30_combout )))

	.dataa(\syif.addr[16]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~30_combout ),
	.cin(gnd),
	.combout(\ramaddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~31 .lut_mask = 16'hBB88;
defparam \ramaddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N2
cycloneive_lcell_comb \ramaddr~32 (
// Equation(s):
// \ramaddr~32_combout  = (temp_dmemWEN1 & (temp_aluResult_19)) # (!temp_dmemWEN1 & ((temp_dmemREN1 & (temp_aluResult_19)) # (!temp_dmemREN1 & ((pccount_19)))))

	.dataa(\CPU|DP|EXMEM|temp_aluResult [19]),
	.datab(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datac(\CPU|DP|PC|pccount [19]),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~32 .lut_mask = 16'hAAB8;
defparam \ramaddr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N20
cycloneive_lcell_comb \ramaddr~33 (
// Equation(s):
// \ramaddr~33_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~32_combout )))

	.dataa(\syif.addr[19]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~32_combout ),
	.cin(gnd),
	.combout(\ramaddr~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~33 .lut_mask = 16'hBB88;
defparam \ramaddr~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N12
cycloneive_lcell_comb \ramaddr~34 (
// Equation(s):
// \ramaddr~34_combout  = (temp_dmemWEN1 & (temp_aluResult_18)) # (!temp_dmemWEN1 & ((temp_dmemREN1 & (temp_aluResult_18)) # (!temp_dmemREN1 & ((pccount_18)))))

	.dataa(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datab(\CPU|DP|EXMEM|temp_aluResult [18]),
	.datac(\CPU|DP|PC|pccount [18]),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~34 .lut_mask = 16'hCCD8;
defparam \ramaddr~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N30
cycloneive_lcell_comb \ramaddr~35 (
// Equation(s):
// \ramaddr~35_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~34_combout )))

	.dataa(gnd),
	.datab(\syif.addr[18]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~34_combout ),
	.cin(gnd),
	.combout(\ramaddr~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~35 .lut_mask = 16'hCFC0;
defparam \ramaddr~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N18
cycloneive_lcell_comb \ramaddr~36 (
// Equation(s):
// \ramaddr~36_combout  = (temp_dmemWEN1 & (temp_aluResult_20)) # (!temp_dmemWEN1 & ((temp_dmemREN1 & (temp_aluResult_20)) # (!temp_dmemREN1 & ((pccount_20)))))

	.dataa(\CPU|DP|EXMEM|temp_aluResult [20]),
	.datab(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datac(\CPU|DP|PC|pccount [20]),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~36 .lut_mask = 16'hAAB8;
defparam \ramaddr~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N30
cycloneive_lcell_comb \ramaddr~37 (
// Equation(s):
// \ramaddr~37_combout  = (temp_dmemREN1 & (temp_aluResult_21)) # (!temp_dmemREN1 & ((temp_dmemWEN1 & (temp_aluResult_21)) # (!temp_dmemWEN1 & ((pccount_21)))))

	.dataa(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datab(\CPU|DP|EXMEM|temp_aluResult [21]),
	.datac(\CPU|DP|PC|pccount [21]),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~37 .lut_mask = 16'hCCD8;
defparam \ramaddr~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N2
cycloneive_lcell_comb \ramaddr~38 (
// Equation(s):
// \ramaddr~38_combout  = (temp_dmemWEN1 & (((temp_aluResult_23)))) # (!temp_dmemWEN1 & ((temp_dmemREN1 & ((temp_aluResult_23))) # (!temp_dmemREN1 & (pccount_23))))

	.dataa(\CPU|DP|PC|pccount [23]),
	.datab(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datac(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datad(\CPU|DP|EXMEM|temp_aluResult [23]),
	.cin(gnd),
	.combout(\ramaddr~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~38 .lut_mask = 16'hFE02;
defparam \ramaddr~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N14
cycloneive_lcell_comb \ramaddr~39 (
// Equation(s):
// \ramaddr~39_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[23]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~38_combout )))

	.dataa(\syif.addr[23]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~38_combout ),
	.cin(gnd),
	.combout(\ramaddr~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~39 .lut_mask = 16'hAFA0;
defparam \ramaddr~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N28
cycloneive_lcell_comb \ramaddr~40 (
// Equation(s):
// \ramaddr~40_combout  = (temp_dmemREN1 & (temp_aluResult_22)) # (!temp_dmemREN1 & ((temp_dmemWEN1 & (temp_aluResult_22)) # (!temp_dmemWEN1 & ((pccount_22)))))

	.dataa(\CPU|DP|EXMEM|temp_aluResult [22]),
	.datab(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datac(\CPU|DP|PC|pccount [22]),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~40 .lut_mask = 16'hAAB8;
defparam \ramaddr~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N22
cycloneive_lcell_comb \ramaddr~41 (
// Equation(s):
// \ramaddr~41_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[22]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~40_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[22]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~40_combout ),
	.cin(gnd),
	.combout(\ramaddr~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~41 .lut_mask = 16'hDD88;
defparam \ramaddr~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N2
cycloneive_lcell_comb \ramaddr~42 (
// Equation(s):
// \ramaddr~42_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[25]~input_o )) # (!\syif.tbCTRL~input_o  & (((temp_dmemWEN1) # (temp_dmemREN1))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[25]~input_o ),
	.datac(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~42 .lut_mask = 16'hDDD8;
defparam \ramaddr~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N18
cycloneive_lcell_comb \ramaddr~43 (
// Equation(s):
// \ramaddr~43_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~42_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~42_combout  & ((temp_aluResult_25))) # (!\ramaddr~42_combout  & (pccount_25))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PC|pccount [25]),
	.datac(\CPU|DP|EXMEM|temp_aluResult [25]),
	.datad(\ramaddr~42_combout ),
	.cin(gnd),
	.combout(\ramaddr~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~43 .lut_mask = 16'hFA44;
defparam \ramaddr~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N20
cycloneive_lcell_comb \ramaddr~44 (
// Equation(s):
// \ramaddr~44_combout  = (temp_dmemWEN1 & (temp_aluResult_24)) # (!temp_dmemWEN1 & ((temp_dmemREN1 & (temp_aluResult_24)) # (!temp_dmemREN1 & ((pccount_24)))))

	.dataa(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datab(\CPU|DP|EXMEM|temp_aluResult [24]),
	.datac(\CPU|DP|PC|pccount [24]),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~44 .lut_mask = 16'hCCD8;
defparam \ramaddr~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N24
cycloneive_lcell_comb \ramaddr~45 (
// Equation(s):
// \ramaddr~45_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~44_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[24]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~44_combout ),
	.cin(gnd),
	.combout(\ramaddr~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~45 .lut_mask = 16'hDD88;
defparam \ramaddr~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N8
cycloneive_lcell_comb \ramaddr~46 (
// Equation(s):
// \ramaddr~46_combout  = (temp_dmemWEN1 & (((temp_aluResult_26)))) # (!temp_dmemWEN1 & ((temp_dmemREN1 & ((temp_aluResult_26))) # (!temp_dmemREN1 & (pccount_26))))

	.dataa(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datab(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datac(\CPU|DP|PC|pccount [26]),
	.datad(\CPU|DP|EXMEM|temp_aluResult [26]),
	.cin(gnd),
	.combout(\ramaddr~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~46 .lut_mask = 16'hFE10;
defparam \ramaddr~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N28
cycloneive_lcell_comb \ramaddr~47 (
// Equation(s):
// \ramaddr~47_combout  = (temp_dmemWEN1 & (temp_aluResult_27)) # (!temp_dmemWEN1 & ((temp_dmemREN1 & (temp_aluResult_27)) # (!temp_dmemREN1 & ((pccount_27)))))

	.dataa(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datab(\CPU|DP|EXMEM|temp_aluResult [27]),
	.datac(\CPU|DP|PC|pccount [27]),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~47 .lut_mask = 16'hCCD8;
defparam \ramaddr~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N0
cycloneive_lcell_comb \ramaddr~48 (
// Equation(s):
// \ramaddr~48_combout  = (temp_dmemWEN1 & (temp_aluResult_29)) # (!temp_dmemWEN1 & ((temp_dmemREN1 & (temp_aluResult_29)) # (!temp_dmemREN1 & ((pccount_29)))))

	.dataa(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datab(\CPU|DP|EXMEM|temp_aluResult [29]),
	.datac(\CPU|DP|PC|pccount [29]),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~48 .lut_mask = 16'hCCD8;
defparam \ramaddr~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N6
cycloneive_lcell_comb \ramaddr~49 (
// Equation(s):
// \ramaddr~49_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[29]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~48_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[29]~input_o ),
	.datad(\ramaddr~48_combout ),
	.cin(gnd),
	.combout(\ramaddr~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~49 .lut_mask = 16'hF3C0;
defparam \ramaddr~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N0
cycloneive_lcell_comb \ramaddr~50 (
// Equation(s):
// \ramaddr~50_combout  = (temp_dmemWEN1 & (temp_aluResult_28)) # (!temp_dmemWEN1 & ((temp_dmemREN1 & (temp_aluResult_28)) # (!temp_dmemREN1 & ((pccount_28)))))

	.dataa(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datab(\CPU|DP|EXMEM|temp_aluResult [28]),
	.datac(\CPU|DP|PC|pccount [28]),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~50 .lut_mask = 16'hCCD8;
defparam \ramaddr~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N12
cycloneive_lcell_comb \ramaddr~51 (
// Equation(s):
// \ramaddr~51_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[28]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~50_combout )))

	.dataa(\syif.addr[28]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~50_combout ),
	.cin(gnd),
	.combout(\ramaddr~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~51 .lut_mask = 16'hBB88;
defparam \ramaddr~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N28
cycloneive_lcell_comb \ramaddr~52 (
// Equation(s):
// \ramaddr~52_combout  = (temp_dmemREN1 & (temp_aluResult_31)) # (!temp_dmemREN1 & ((temp_dmemWEN1 & (temp_aluResult_31)) # (!temp_dmemWEN1 & ((pccount_31)))))

	.dataa(\CPU|DP|EXMEM|temp_aluResult [31]),
	.datab(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datac(\CPU|DP|PC|pccount [31]),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~52 .lut_mask = 16'hAAB8;
defparam \ramaddr~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N30
cycloneive_lcell_comb \ramaddr~53 (
// Equation(s):
// \ramaddr~53_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~52_combout )))

	.dataa(gnd),
	.datab(\syif.addr[31]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~52_combout ),
	.cin(gnd),
	.combout(\ramaddr~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~53 .lut_mask = 16'hCFC0;
defparam \ramaddr~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N8
cycloneive_lcell_comb \ramaddr~54 (
// Equation(s):
// \ramaddr~54_combout  = (temp_dmemWEN1 & (temp_aluResult_30)) # (!temp_dmemWEN1 & ((temp_dmemREN1 & (temp_aluResult_30)) # (!temp_dmemREN1 & ((pccount_30)))))

	.dataa(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datab(\CPU|DP|EXMEM|temp_aluResult [30]),
	.datac(\CPU|DP|PC|pccount [30]),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~54 .lut_mask = 16'hCCD8;
defparam \ramaddr~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N28
cycloneive_lcell_comb \ramaddr~55 (
// Equation(s):
// \ramaddr~55_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[30]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~54_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[30]~input_o ),
	.datad(\ramaddr~54_combout ),
	.cin(gnd),
	.combout(\ramaddr~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~55 .lut_mask = 16'hF5A0;
defparam \ramaddr~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y72_N11
dffeas CPUCLK(
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\CPUCLK~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\CPUCLK~q ),
	.prn(vcc));
// synopsys translate_off
defparam CPUCLK.is_wysiwyg = "true";
defparam CPUCLK.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N14
cycloneive_lcell_comb \ramWEN~0 (
// Equation(s):
// \ramWEN~0_combout  = (\syif.tbCTRL~input_o  & (((\syif.WEN~input_o )))) # (!\syif.tbCTRL~input_o  & (temp_dmemWEN1 & ((!temp_dmemREN1))))

	.dataa(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datab(\syif.WEN~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramWEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramWEN~0 .lut_mask = 16'hC0CA;
defparam \ramWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N22
cycloneive_lcell_comb \ramWEN~1 (
// Equation(s):
// \ramWEN~1_combout  = (!\syif.tbCTRL~input_o  & (temp_dmemWEN1 & !temp_dmemREN1))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.datad(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.cin(gnd),
	.combout(\ramWEN~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramWEN~1 .lut_mask = 16'h0030;
defparam \ramWEN~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N8
cycloneive_lcell_comb \ramstore~0 (
// Equation(s):
// \ramstore~0_combout  = (\syif.store[0]~input_o  & ((\syif.tbCTRL~input_o ) # ((\ramWEN~1_combout  & temp_rdat2_0)))) # (!\syif.store[0]~input_o  & (((\ramWEN~1_combout  & temp_rdat2_0))))

	.dataa(\syif.store[0]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramWEN~1_combout ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [0]),
	.cin(gnd),
	.combout(\ramstore~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~0 .lut_mask = 16'hF888;
defparam \ramstore~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N4
cycloneive_lcell_comb \ramaddr~56 (
// Equation(s):
// \ramaddr~56_combout  = (\syif.tbCTRL~input_o  & ((\syif.addr[2]~input_o ))) # (!\syif.tbCTRL~input_o  & (\ramaddr~2_combout ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\ramaddr~2_combout ),
	.datac(gnd),
	.datad(\syif.addr[2]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~56 .lut_mask = 16'hEE44;
defparam \ramaddr~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N8
cycloneive_lcell_comb \ramaddr~57 (
// Equation(s):
// \ramaddr~57_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[3]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~3_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[3]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~3_combout ),
	.cin(gnd),
	.combout(\ramaddr~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~57 .lut_mask = 16'hDD88;
defparam \ramaddr~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N30
cycloneive_lcell_comb \ramaddr~58 (
// Equation(s):
// \ramaddr~58_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~1_combout )))

	.dataa(gnd),
	.datab(\syif.addr[0]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~1_combout ),
	.cin(gnd),
	.combout(\ramaddr~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~58 .lut_mask = 16'hCFC0;
defparam \ramaddr~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N0
cycloneive_lcell_comb \ramaddr~59 (
// Equation(s):
// \ramaddr~59_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[1]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~0_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[1]~input_o ),
	.datac(\ramaddr~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramaddr~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~59 .lut_mask = 16'hD8D8;
defparam \ramaddr~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N4
cycloneive_lcell_comb \ramaddr~60 (
// Equation(s):
// \ramaddr~60_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[21]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~37_combout )))

	.dataa(gnd),
	.datab(\syif.addr[21]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~37_combout ),
	.cin(gnd),
	.combout(\ramaddr~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~60 .lut_mask = 16'hCFC0;
defparam \ramaddr~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N16
cycloneive_lcell_comb \ramaddr~61 (
// Equation(s):
// \ramaddr~61_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~36_combout )))

	.dataa(gnd),
	.datab(\syif.addr[20]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~36_combout ),
	.cin(gnd),
	.combout(\ramaddr~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~61 .lut_mask = 16'hCFC0;
defparam \ramaddr~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N30
cycloneive_lcell_comb \ramaddr~62 (
// Equation(s):
// \ramaddr~62_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~47_combout )))

	.dataa(\syif.addr[27]~input_o ),
	.datab(\ramaddr~47_combout ),
	.datac(gnd),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~62 .lut_mask = 16'hAACC;
defparam \ramaddr~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N16
cycloneive_lcell_comb \ramaddr~63 (
// Equation(s):
// \ramaddr~63_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[26]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~46_combout )))

	.dataa(\syif.addr[26]~input_o ),
	.datab(gnd),
	.datac(\ramaddr~46_combout ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~63 .lut_mask = 16'hAAF0;
defparam \ramaddr~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N30
cycloneive_lcell_comb \ramstore~1 (
// Equation(s):
// \ramstore~1_combout  = (\ramWEN~1_combout  & ((temp_rdat2_1) # ((\syif.tbCTRL~input_o  & \syif.store[1]~input_o )))) # (!\ramWEN~1_combout  & (\syif.tbCTRL~input_o  & ((\syif.store[1]~input_o ))))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|temp_rdat2 [1]),
	.datad(\syif.store[1]~input_o ),
	.cin(gnd),
	.combout(\ramstore~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~1 .lut_mask = 16'hECA0;
defparam \ramstore~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N20
cycloneive_lcell_comb \ramstore~2 (
// Equation(s):
// \ramstore~2_combout  = (\ramWEN~1_combout  & ((temp_rdat2_2) # ((\syif.store[2]~input_o  & \syif.tbCTRL~input_o )))) # (!\ramWEN~1_combout  & (\syif.store[2]~input_o  & (\syif.tbCTRL~input_o )))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.store[2]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [2]),
	.cin(gnd),
	.combout(\ramstore~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~2 .lut_mask = 16'hEAC0;
defparam \ramstore~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N12
cycloneive_lcell_comb \ramstore~3 (
// Equation(s):
// \ramstore~3_combout  = (\syif.store[3]~input_o  & ((\syif.tbCTRL~input_o ) # ((\ramWEN~1_combout  & temp_rdat2_3)))) # (!\syif.store[3]~input_o  & (((\ramWEN~1_combout  & temp_rdat2_3))))

	.dataa(\syif.store[3]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramWEN~1_combout ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [3]),
	.cin(gnd),
	.combout(\ramstore~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~3 .lut_mask = 16'hF888;
defparam \ramstore~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N6
cycloneive_lcell_comb \ramstore~4 (
// Equation(s):
// \ramstore~4_combout  = (\ramWEN~1_combout  & ((temp_rdat2_4) # ((\syif.tbCTRL~input_o  & \syif.store[4]~input_o )))) # (!\ramWEN~1_combout  & (((\syif.tbCTRL~input_o  & \syif.store[4]~input_o ))))

	.dataa(\ramWEN~1_combout ),
	.datab(\CPU|DP|EXMEM|temp_rdat2 [4]),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\syif.store[4]~input_o ),
	.cin(gnd),
	.combout(\ramstore~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~4 .lut_mask = 16'hF888;
defparam \ramstore~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N18
cycloneive_lcell_comb \ramstore~5 (
// Equation(s):
// \ramstore~5_combout  = (temp_rdat2_5 & ((\ramWEN~1_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[5]~input_o )))) # (!temp_rdat2_5 & (\syif.tbCTRL~input_o  & ((\syif.store[5]~input_o ))))

	.dataa(\CPU|DP|EXMEM|temp_rdat2 [5]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramWEN~1_combout ),
	.datad(\syif.store[5]~input_o ),
	.cin(gnd),
	.combout(\ramstore~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~5 .lut_mask = 16'hECA0;
defparam \ramstore~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N28
cycloneive_lcell_comb \ramstore~6 (
// Equation(s):
// \ramstore~6_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[6]~input_o ) # ((temp_rdat2_6 & \ramWEN~1_combout )))) # (!\syif.tbCTRL~input_o  & (temp_rdat2_6 & (\ramWEN~1_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|temp_rdat2 [6]),
	.datac(\ramWEN~1_combout ),
	.datad(\syif.store[6]~input_o ),
	.cin(gnd),
	.combout(\ramstore~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~6 .lut_mask = 16'hEAC0;
defparam \ramstore~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N0
cycloneive_lcell_comb \ramstore~7 (
// Equation(s):
// \ramstore~7_combout  = (temp_rdat2_7 & ((\ramWEN~1_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[7]~input_o )))) # (!temp_rdat2_7 & (\syif.tbCTRL~input_o  & ((\syif.store[7]~input_o ))))

	.dataa(\CPU|DP|EXMEM|temp_rdat2 [7]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramWEN~1_combout ),
	.datad(\syif.store[7]~input_o ),
	.cin(gnd),
	.combout(\ramstore~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~7 .lut_mask = 16'hECA0;
defparam \ramstore~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N2
cycloneive_lcell_comb \ramstore~8 (
// Equation(s):
// \ramstore~8_combout  = (\syif.store[8]~input_o  & ((\syif.tbCTRL~input_o ) # ((\ramWEN~1_combout  & temp_rdat2_8)))) # (!\syif.store[8]~input_o  & (((\ramWEN~1_combout  & temp_rdat2_8))))

	.dataa(\syif.store[8]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramWEN~1_combout ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [8]),
	.cin(gnd),
	.combout(\ramstore~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~8 .lut_mask = 16'hF888;
defparam \ramstore~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N2
cycloneive_lcell_comb \ramstore~9 (
// Equation(s):
// \ramstore~9_combout  = (\ramWEN~1_combout  & ((temp_rdat2_9) # ((\syif.store[9]~input_o  & \syif.tbCTRL~input_o )))) # (!\ramWEN~1_combout  & (\syif.store[9]~input_o  & (\syif.tbCTRL~input_o )))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.store[9]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [9]),
	.cin(gnd),
	.combout(\ramstore~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~9 .lut_mask = 16'hEAC0;
defparam \ramstore~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N28
cycloneive_lcell_comb \ramstore~10 (
// Equation(s):
// \ramstore~10_combout  = (\syif.store[10]~input_o  & ((\syif.tbCTRL~input_o ) # ((\ramWEN~1_combout  & temp_rdat2_10)))) # (!\syif.store[10]~input_o  & (((\ramWEN~1_combout  & temp_rdat2_10))))

	.dataa(\syif.store[10]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramWEN~1_combout ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [10]),
	.cin(gnd),
	.combout(\ramstore~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~10 .lut_mask = 16'hF888;
defparam \ramstore~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N10
cycloneive_lcell_comb \ramstore~11 (
// Equation(s):
// \ramstore~11_combout  = (\syif.store[11]~input_o  & ((\syif.tbCTRL~input_o ) # ((temp_rdat2_11 & \ramWEN~1_combout )))) # (!\syif.store[11]~input_o  & (temp_rdat2_11 & (\ramWEN~1_combout )))

	.dataa(\syif.store[11]~input_o ),
	.datab(\CPU|DP|EXMEM|temp_rdat2 [11]),
	.datac(\ramWEN~1_combout ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~11 .lut_mask = 16'hEAC0;
defparam \ramstore~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N20
cycloneive_lcell_comb \ramstore~12 (
// Equation(s):
// \ramstore~12_combout  = (temp_rdat2_12 & ((\ramWEN~1_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[12]~input_o )))) # (!temp_rdat2_12 & (\syif.tbCTRL~input_o  & ((\syif.store[12]~input_o ))))

	.dataa(\CPU|DP|EXMEM|temp_rdat2 [12]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramWEN~1_combout ),
	.datad(\syif.store[12]~input_o ),
	.cin(gnd),
	.combout(\ramstore~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~12 .lut_mask = 16'hECA0;
defparam \ramstore~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N6
cycloneive_lcell_comb \ramstore~13 (
// Equation(s):
// \ramstore~13_combout  = (temp_rdat2_13 & ((\ramWEN~1_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[13]~input_o )))) # (!temp_rdat2_13 & (\syif.tbCTRL~input_o  & ((\syif.store[13]~input_o ))))

	.dataa(\CPU|DP|EXMEM|temp_rdat2 [13]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramWEN~1_combout ),
	.datad(\syif.store[13]~input_o ),
	.cin(gnd),
	.combout(\ramstore~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~13 .lut_mask = 16'hECA0;
defparam \ramstore~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N4
cycloneive_lcell_comb \ramstore~14 (
// Equation(s):
// \ramstore~14_combout  = (\ramWEN~1_combout  & ((temp_rdat2_14) # ((\syif.store[14]~input_o  & \syif.tbCTRL~input_o )))) # (!\ramWEN~1_combout  & (\syif.store[14]~input_o  & ((\syif.tbCTRL~input_o ))))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.store[14]~input_o ),
	.datac(\CPU|DP|EXMEM|temp_rdat2 [14]),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~14 .lut_mask = 16'hECA0;
defparam \ramstore~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N26
cycloneive_lcell_comb \ramstore~15 (
// Equation(s):
// \ramstore~15_combout  = (\syif.store[15]~input_o  & ((\syif.tbCTRL~input_o ) # ((temp_rdat2_15 & \ramWEN~1_combout )))) # (!\syif.store[15]~input_o  & (temp_rdat2_15 & (\ramWEN~1_combout )))

	.dataa(\syif.store[15]~input_o ),
	.datab(\CPU|DP|EXMEM|temp_rdat2 [15]),
	.datac(\ramWEN~1_combout ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~15 .lut_mask = 16'hEAC0;
defparam \ramstore~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N24
cycloneive_lcell_comb \ramstore~16 (
// Equation(s):
// \ramstore~16_combout  = (\ramWEN~1_combout  & ((temp_rdat2_16) # ((\syif.tbCTRL~input_o  & \syif.store[16]~input_o )))) # (!\ramWEN~1_combout  & (\syif.tbCTRL~input_o  & (\syif.store[16]~input_o )))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[16]~input_o ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [16]),
	.cin(gnd),
	.combout(\ramstore~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~16 .lut_mask = 16'hEAC0;
defparam \ramstore~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N18
cycloneive_lcell_comb \ramstore~17 (
// Equation(s):
// \ramstore~17_combout  = (\ramWEN~1_combout  & ((temp_rdat2_17) # ((\syif.tbCTRL~input_o  & \syif.store[17]~input_o )))) # (!\ramWEN~1_combout  & (\syif.tbCTRL~input_o  & (\syif.store[17]~input_o )))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[17]~input_o ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [17]),
	.cin(gnd),
	.combout(\ramstore~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~17 .lut_mask = 16'hEAC0;
defparam \ramstore~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N24
cycloneive_lcell_comb \ramstore~18 (
// Equation(s):
// \ramstore~18_combout  = (temp_rdat2_18 & ((\ramWEN~1_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[18]~input_o )))) # (!temp_rdat2_18 & (\syif.tbCTRL~input_o  & ((\syif.store[18]~input_o ))))

	.dataa(\CPU|DP|EXMEM|temp_rdat2 [18]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramWEN~1_combout ),
	.datad(\syif.store[18]~input_o ),
	.cin(gnd),
	.combout(\ramstore~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~18 .lut_mask = 16'hECA0;
defparam \ramstore~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N0
cycloneive_lcell_comb \ramstore~19 (
// Equation(s):
// \ramstore~19_combout  = (\ramWEN~1_combout  & ((temp_rdat2_19) # ((\syif.store[19]~input_o  & \syif.tbCTRL~input_o )))) # (!\ramWEN~1_combout  & (\syif.store[19]~input_o  & (\syif.tbCTRL~input_o )))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.store[19]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [19]),
	.cin(gnd),
	.combout(\ramstore~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~19 .lut_mask = 16'hEAC0;
defparam \ramstore~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N18
cycloneive_lcell_comb \ramstore~20 (
// Equation(s):
// \ramstore~20_combout  = (\ramWEN~1_combout  & ((temp_rdat2_20) # ((\syif.store[20]~input_o  & \syif.tbCTRL~input_o )))) # (!\ramWEN~1_combout  & (\syif.store[20]~input_o  & (\syif.tbCTRL~input_o )))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.store[20]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [20]),
	.cin(gnd),
	.combout(\ramstore~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~20 .lut_mask = 16'hEAC0;
defparam \ramstore~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N24
cycloneive_lcell_comb \ramstore~21 (
// Equation(s):
// \ramstore~21_combout  = (\ramWEN~1_combout  & ((temp_rdat2_21) # ((\syif.store[21]~input_o  & \syif.tbCTRL~input_o )))) # (!\ramWEN~1_combout  & (\syif.store[21]~input_o  & (\syif.tbCTRL~input_o )))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.store[21]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [21]),
	.cin(gnd),
	.combout(\ramstore~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~21 .lut_mask = 16'hEAC0;
defparam \ramstore~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N26
cycloneive_lcell_comb \ramstore~22 (
// Equation(s):
// \ramstore~22_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[22]~input_o ) # ((\ramWEN~1_combout  & temp_rdat2_22)))) # (!\syif.tbCTRL~input_o  & (((\ramWEN~1_combout  & temp_rdat2_22))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[22]~input_o ),
	.datac(\ramWEN~1_combout ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [22]),
	.cin(gnd),
	.combout(\ramstore~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~22 .lut_mask = 16'hF888;
defparam \ramstore~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N22
cycloneive_lcell_comb \ramstore~23 (
// Equation(s):
// \ramstore~23_combout  = (\syif.store[23]~input_o  & ((\syif.tbCTRL~input_o ) # ((temp_rdat2_23 & \ramWEN~1_combout )))) # (!\syif.store[23]~input_o  & (temp_rdat2_23 & (\ramWEN~1_combout )))

	.dataa(\syif.store[23]~input_o ),
	.datab(\CPU|DP|EXMEM|temp_rdat2 [23]),
	.datac(\ramWEN~1_combout ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~23 .lut_mask = 16'hEAC0;
defparam \ramstore~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N22
cycloneive_lcell_comb \ramstore~24 (
// Equation(s):
// \ramstore~24_combout  = (\ramWEN~1_combout  & ((temp_rdat2_24) # ((\syif.store[24]~input_o  & \syif.tbCTRL~input_o )))) # (!\ramWEN~1_combout  & (\syif.store[24]~input_o  & (\syif.tbCTRL~input_o )))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.store[24]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [24]),
	.cin(gnd),
	.combout(\ramstore~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~24 .lut_mask = 16'hEAC0;
defparam \ramstore~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N22
cycloneive_lcell_comb \ramstore~25 (
// Equation(s):
// \ramstore~25_combout  = (\syif.store[25]~input_o  & ((\syif.tbCTRL~input_o ) # ((temp_rdat2_25 & \ramWEN~1_combout )))) # (!\syif.store[25]~input_o  & (((temp_rdat2_25 & \ramWEN~1_combout ))))

	.dataa(\syif.store[25]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|temp_rdat2 [25]),
	.datad(\ramWEN~1_combout ),
	.cin(gnd),
	.combout(\ramstore~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~25 .lut_mask = 16'hF888;
defparam \ramstore~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N16
cycloneive_lcell_comb \ramstore~26 (
// Equation(s):
// \ramstore~26_combout  = (\ramWEN~1_combout  & ((temp_rdat2_26) # ((\syif.tbCTRL~input_o  & \syif.store[26]~input_o )))) # (!\ramWEN~1_combout  & (((\syif.tbCTRL~input_o  & \syif.store[26]~input_o ))))

	.dataa(\ramWEN~1_combout ),
	.datab(\CPU|DP|EXMEM|temp_rdat2 [26]),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\syif.store[26]~input_o ),
	.cin(gnd),
	.combout(\ramstore~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~26 .lut_mask = 16'hF888;
defparam \ramstore~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N10
cycloneive_lcell_comb \ramstore~27 (
// Equation(s):
// \ramstore~27_combout  = (\ramWEN~1_combout  & ((temp_rdat2_27) # ((\syif.tbCTRL~input_o  & \syif.store[27]~input_o )))) # (!\ramWEN~1_combout  & (((\syif.tbCTRL~input_o  & \syif.store[27]~input_o ))))

	.dataa(\ramWEN~1_combout ),
	.datab(\CPU|DP|EXMEM|temp_rdat2 [27]),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\syif.store[27]~input_o ),
	.cin(gnd),
	.combout(\ramstore~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~27 .lut_mask = 16'hF888;
defparam \ramstore~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N22
cycloneive_lcell_comb \ramstore~28 (
// Equation(s):
// \ramstore~28_combout  = (\ramWEN~1_combout  & ((temp_rdat2_28) # ((\syif.store[28]~input_o  & \syif.tbCTRL~input_o )))) # (!\ramWEN~1_combout  & (((\syif.store[28]~input_o  & \syif.tbCTRL~input_o ))))

	.dataa(\ramWEN~1_combout ),
	.datab(\CPU|DP|EXMEM|temp_rdat2 [28]),
	.datac(\syif.store[28]~input_o ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~28 .lut_mask = 16'hF888;
defparam \ramstore~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N12
cycloneive_lcell_comb \ramstore~29 (
// Equation(s):
// \ramstore~29_combout  = (\ramWEN~1_combout  & ((temp_rdat2_29) # ((\syif.store[29]~input_o  & \syif.tbCTRL~input_o )))) # (!\ramWEN~1_combout  & (\syif.store[29]~input_o  & (\syif.tbCTRL~input_o )))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.store[29]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [29]),
	.cin(gnd),
	.combout(\ramstore~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~29 .lut_mask = 16'hEAC0;
defparam \ramstore~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N16
cycloneive_lcell_comb \ramstore~30 (
// Equation(s):
// \ramstore~30_combout  = (\syif.store[30]~input_o  & ((\syif.tbCTRL~input_o ) # ((\ramWEN~1_combout  & temp_rdat2_30)))) # (!\syif.store[30]~input_o  & (((\ramWEN~1_combout  & temp_rdat2_30))))

	.dataa(\syif.store[30]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramWEN~1_combout ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [30]),
	.cin(gnd),
	.combout(\ramstore~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~30 .lut_mask = 16'hF888;
defparam \ramstore~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N26
cycloneive_lcell_comb \ramstore~31 (
// Equation(s):
// \ramstore~31_combout  = (\ramWEN~1_combout  & ((temp_rdat2_31) # ((\syif.store[31]~input_o  & \syif.tbCTRL~input_o )))) # (!\ramWEN~1_combout  & (\syif.store[31]~input_o  & (\syif.tbCTRL~input_o )))

	.dataa(\ramWEN~1_combout ),
	.datab(\syif.store[31]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|temp_rdat2 [31]),
	.cin(gnd),
	.combout(\ramstore~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~31 .lut_mask = 16'hEAC0;
defparam \ramstore~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y72_N1
dffeas \count[3] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y72_N7
dffeas \count[2] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y72_N9
dffeas \count[1] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y72_N19
dffeas \count[0] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N12
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!count[2] & (!count[0] & (!count[1] & !count[3])))

	.dataa(count[2]),
	.datab(count[0]),
	.datac(count[1]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h0001;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N10
cycloneive_lcell_comb \CPUCLK~0 (
// Equation(s):
// \CPUCLK~0_combout  = \CPUCLK~q  $ (\Equal0~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\CPUCLK~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\CPUCLK~0_combout ),
	.cout());
// synopsys translate_off
defparam \CPUCLK~0 .lut_mask = 16'h0FF0;
defparam \CPUCLK~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N6
cycloneive_lcell_comb \ramREN~0 (
// Equation(s):
// \ramREN~0_combout  = (\syif.tbCTRL~input_o  & (\syif.REN~input_o )) # (!\syif.tbCTRL~input_o  & (((temp_dmemREN1) # (!temp_dmemWEN1))))

	.dataa(\syif.REN~input_o ),
	.datab(\CPU|DP|EXMEM|temp_dmemREN~q ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|temp_dmemWEN~q ),
	.cin(gnd),
	.combout(\ramREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramREN~0 .lut_mask = 16'hACAF;
defparam \ramREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N0
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = count[3] $ (((count[2] & (count[1] & count[0]))))

	.dataa(count[2]),
	.datab(count[1]),
	.datac(count[3]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h78F0;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N6
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = count[2] $ (((count[1] & count[0])))

	.dataa(gnd),
	.datab(count[1]),
	.datac(count[2]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h3CF0;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N8
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = count[1] $ (count[0])

	.dataa(gnd),
	.datab(gnd),
	.datac(count[1]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h0FF0;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N18
cycloneive_lcell_comb \count~3 (
// Equation(s):
// \count~3_combout  = (!count[0] & ((count[2]) # ((count[1]) # (count[3]))))

	.dataa(count[2]),
	.datab(count[1]),
	.datac(count[0]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
// synopsys translate_off
defparam \count~3 .lut_mask = 16'h0F0E;
defparam \count~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N8
cycloneive_lcell_comb \ramaddr~25_wirecell (
// Equation(s):
// \ramaddr~25_wirecell_combout  = !\ramaddr~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\ramaddr~25_combout ),
	.cin(gnd),
	.combout(\ramaddr~25_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~25_wirecell .lut_mask = 16'h00FF;
defparam \ramaddr~25_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: JTAG_X1_Y37_N0
cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

// Location: FF_X46_Y40_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y40_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y42_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y40_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .lut_mask = 16'h55AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X45_Y41_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y41_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y41_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y41_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y41_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y40_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datab(gnd),
	.datac(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .lut_mask = 16'hF0AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .lut_mask = 16'hAAB0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .lut_mask = 16'hFFA0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .lut_mask = 16'hA0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .lut_mask = 16'hDF80;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .lut_mask = 16'h040C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .lut_mask = 16'hEE20;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .lut_mask = 16'hAA30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .lut_mask = 16'h0001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .lut_mask = 16'hFAFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .lut_mask = 16'hC001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .lut_mask = 16'h0002;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .lut_mask = 16'h4CCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .lut_mask = 16'h0C0D;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 .lut_mask = 16'hCFC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y40_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .lut_mask = 16'hFF40;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .lut_mask = 16'hF0F1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .lut_mask = 16'h9746;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .lut_mask = 16'h00F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .lut_mask = 16'h192D;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .lut_mask = 16'h0C7C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N8
cycloneive_io_ibuf \syif.WEN~input (
	.i(\syif.WEN ),
	.ibar(gnd),
	.o(\syif.WEN~input_o ));
// synopsys translate_off
defparam \syif.WEN~input .bus_hold = "false";
defparam \syif.WEN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N1
cycloneive_io_ibuf \syif.tbCTRL~input (
	.i(\syif.tbCTRL ),
	.ibar(gnd),
	.o(\syif.tbCTRL~input_o ));
// synopsys translate_off
defparam \syif.tbCTRL~input .bus_hold = "false";
defparam \syif.tbCTRL~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N8
cycloneive_io_ibuf \syif.REN~input (
	.i(\syif.REN ),
	.ibar(gnd),
	.o(\syif.REN~input_o ));
// synopsys translate_off
defparam \syif.REN~input .bus_hold = "false";
defparam \syif.REN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y73_N22
cycloneive_io_ibuf \syif.addr[0]~input (
	.i(\syif.addr [0]),
	.ibar(gnd),
	.o(\syif.addr[0]~input_o ));
// synopsys translate_off
defparam \syif.addr[0]~input .bus_hold = "false";
defparam \syif.addr[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N22
cycloneive_io_ibuf \syif.addr[1]~input (
	.i(\syif.addr [1]),
	.ibar(gnd),
	.o(\syif.addr[1]~input_o ));
// synopsys translate_off
defparam \syif.addr[1]~input .bus_hold = "false";
defparam \syif.addr[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N15
cycloneive_io_ibuf \syif.addr[3]~input (
	.i(\syif.addr [3]),
	.ibar(gnd),
	.o(\syif.addr[3]~input_o ));
// synopsys translate_off
defparam \syif.addr[3]~input .bus_hold = "false";
defparam \syif.addr[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N8
cycloneive_io_ibuf \syif.addr[2]~input (
	.i(\syif.addr [2]),
	.ibar(gnd),
	.o(\syif.addr[2]~input_o ));
// synopsys translate_off
defparam \syif.addr[2]~input .bus_hold = "false";
defparam \syif.addr[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N22
cycloneive_io_ibuf \syif.addr[5]~input (
	.i(\syif.addr [5]),
	.ibar(gnd),
	.o(\syif.addr[5]~input_o ));
// synopsys translate_off
defparam \syif.addr[5]~input .bus_hold = "false";
defparam \syif.addr[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y43_N15
cycloneive_io_ibuf \syif.addr[4]~input (
	.i(\syif.addr [4]),
	.ibar(gnd),
	.o(\syif.addr[4]~input_o ));
// synopsys translate_off
defparam \syif.addr[4]~input .bus_hold = "false";
defparam \syif.addr[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N1
cycloneive_io_ibuf \syif.addr[7]~input (
	.i(\syif.addr [7]),
	.ibar(gnd),
	.o(\syif.addr[7]~input_o ));
// synopsys translate_off
defparam \syif.addr[7]~input .bus_hold = "false";
defparam \syif.addr[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N8
cycloneive_io_ibuf \syif.addr[6]~input (
	.i(\syif.addr [6]),
	.ibar(gnd),
	.o(\syif.addr[6]~input_o ));
// synopsys translate_off
defparam \syif.addr[6]~input .bus_hold = "false";
defparam \syif.addr[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N22
cycloneive_io_ibuf \syif.addr[9]~input (
	.i(\syif.addr [9]),
	.ibar(gnd),
	.o(\syif.addr[9]~input_o ));
// synopsys translate_off
defparam \syif.addr[9]~input .bus_hold = "false";
defparam \syif.addr[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N22
cycloneive_io_ibuf \syif.addr[8]~input (
	.i(\syif.addr [8]),
	.ibar(gnd),
	.o(\syif.addr[8]~input_o ));
// synopsys translate_off
defparam \syif.addr[8]~input .bus_hold = "false";
defparam \syif.addr[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y44_N8
cycloneive_io_ibuf \syif.addr[11]~input (
	.i(\syif.addr [11]),
	.ibar(gnd),
	.o(\syif.addr[11]~input_o ));
// synopsys translate_off
defparam \syif.addr[11]~input .bus_hold = "false";
defparam \syif.addr[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y42_N15
cycloneive_io_ibuf \syif.addr[10]~input (
	.i(\syif.addr [10]),
	.ibar(gnd),
	.o(\syif.addr[10]~input_o ));
// synopsys translate_off
defparam \syif.addr[10]~input .bus_hold = "false";
defparam \syif.addr[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y0_N15
cycloneive_io_ibuf \syif.addr[13]~input (
	.i(\syif.addr [13]),
	.ibar(gnd),
	.o(\syif.addr[13]~input_o ));
// synopsys translate_off
defparam \syif.addr[13]~input .bus_hold = "false";
defparam \syif.addr[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N1
cycloneive_io_ibuf \syif.addr[12]~input (
	.i(\syif.addr [12]),
	.ibar(gnd),
	.o(\syif.addr[12]~input_o ));
// synopsys translate_off
defparam \syif.addr[12]~input .bus_hold = "false";
defparam \syif.addr[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N15
cycloneive_io_ibuf \syif.addr[15]~input (
	.i(\syif.addr [15]),
	.ibar(gnd),
	.o(\syif.addr[15]~input_o ));
// synopsys translate_off
defparam \syif.addr[15]~input .bus_hold = "false";
defparam \syif.addr[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N1
cycloneive_io_ibuf \syif.addr[14]~input (
	.i(\syif.addr [14]),
	.ibar(gnd),
	.o(\syif.addr[14]~input_o ));
// synopsys translate_off
defparam \syif.addr[14]~input .bus_hold = "false";
defparam \syif.addr[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N22
cycloneive_io_ibuf \syif.addr[17]~input (
	.i(\syif.addr [17]),
	.ibar(gnd),
	.o(\syif.addr[17]~input_o ));
// synopsys translate_off
defparam \syif.addr[17]~input .bus_hold = "false";
defparam \syif.addr[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N22
cycloneive_io_ibuf \syif.addr[16]~input (
	.i(\syif.addr [16]),
	.ibar(gnd),
	.o(\syif.addr[16]~input_o ));
// synopsys translate_off
defparam \syif.addr[16]~input .bus_hold = "false";
defparam \syif.addr[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N1
cycloneive_io_ibuf \syif.addr[19]~input (
	.i(\syif.addr [19]),
	.ibar(gnd),
	.o(\syif.addr[19]~input_o ));
// synopsys translate_off
defparam \syif.addr[19]~input .bus_hold = "false";
defparam \syif.addr[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N15
cycloneive_io_ibuf \syif.addr[18]~input (
	.i(\syif.addr [18]),
	.ibar(gnd),
	.o(\syif.addr[18]~input_o ));
// synopsys translate_off
defparam \syif.addr[18]~input .bus_hold = "false";
defparam \syif.addr[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N8
cycloneive_io_ibuf \syif.addr[21]~input (
	.i(\syif.addr [21]),
	.ibar(gnd),
	.o(\syif.addr[21]~input_o ));
// synopsys translate_off
defparam \syif.addr[21]~input .bus_hold = "false";
defparam \syif.addr[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N15
cycloneive_io_ibuf \syif.addr[20]~input (
	.i(\syif.addr [20]),
	.ibar(gnd),
	.o(\syif.addr[20]~input_o ));
// synopsys translate_off
defparam \syif.addr[20]~input .bus_hold = "false";
defparam \syif.addr[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N8
cycloneive_io_ibuf \syif.addr[23]~input (
	.i(\syif.addr [23]),
	.ibar(gnd),
	.o(\syif.addr[23]~input_o ));
// synopsys translate_off
defparam \syif.addr[23]~input .bus_hold = "false";
defparam \syif.addr[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N22
cycloneive_io_ibuf \syif.addr[22]~input (
	.i(\syif.addr [22]),
	.ibar(gnd),
	.o(\syif.addr[22]~input_o ));
// synopsys translate_off
defparam \syif.addr[22]~input .bus_hold = "false";
defparam \syif.addr[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y44_N8
cycloneive_io_ibuf \syif.addr[25]~input (
	.i(\syif.addr [25]),
	.ibar(gnd),
	.o(\syif.addr[25]~input_o ));
// synopsys translate_off
defparam \syif.addr[25]~input .bus_hold = "false";
defparam \syif.addr[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y44_N1
cycloneive_io_ibuf \syif.addr[24]~input (
	.i(\syif.addr [24]),
	.ibar(gnd),
	.o(\syif.addr[24]~input_o ));
// synopsys translate_off
defparam \syif.addr[24]~input .bus_hold = "false";
defparam \syif.addr[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N8
cycloneive_io_ibuf \syif.addr[27]~input (
	.i(\syif.addr [27]),
	.ibar(gnd),
	.o(\syif.addr[27]~input_o ));
// synopsys translate_off
defparam \syif.addr[27]~input .bus_hold = "false";
defparam \syif.addr[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N15
cycloneive_io_ibuf \syif.addr[26]~input (
	.i(\syif.addr [26]),
	.ibar(gnd),
	.o(\syif.addr[26]~input_o ));
// synopsys translate_off
defparam \syif.addr[26]~input .bus_hold = "false";
defparam \syif.addr[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y43_N8
cycloneive_io_ibuf \syif.addr[29]~input (
	.i(\syif.addr [29]),
	.ibar(gnd),
	.o(\syif.addr[29]~input_o ));
// synopsys translate_off
defparam \syif.addr[29]~input .bus_hold = "false";
defparam \syif.addr[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N1
cycloneive_io_ibuf \syif.addr[28]~input (
	.i(\syif.addr [28]),
	.ibar(gnd),
	.o(\syif.addr[28]~input_o ));
// synopsys translate_off
defparam \syif.addr[28]~input .bus_hold = "false";
defparam \syif.addr[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N1
cycloneive_io_ibuf \syif.addr[31]~input (
	.i(\syif.addr [31]),
	.ibar(gnd),
	.o(\syif.addr[31]~input_o ));
// synopsys translate_off
defparam \syif.addr[31]~input .bus_hold = "false";
defparam \syif.addr[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N15
cycloneive_io_ibuf \syif.addr[30]~input (
	.i(\syif.addr [30]),
	.ibar(gnd),
	.o(\syif.addr[30]~input_o ));
// synopsys translate_off
defparam \syif.addr[30]~input .bus_hold = "false";
defparam \syif.addr[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N15
cycloneive_io_ibuf \nRST~input (
	.i(nRST),
	.ibar(gnd),
	.o(\nRST~input_o ));
// synopsys translate_off
defparam \nRST~input .bus_hold = "false";
defparam \nRST~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N8
cycloneive_io_ibuf \CLK~input (
	.i(CLK),
	.ibar(gnd),
	.o(\CLK~input_o ));
// synopsys translate_off
defparam \CLK~input .bus_hold = "false";
defparam \CLK~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N1
cycloneive_io_ibuf \syif.store[0]~input (
	.i(\syif.store [0]),
	.ibar(gnd),
	.o(\syif.store[0]~input_o ));
// synopsys translate_off
defparam \syif.store[0]~input .bus_hold = "false";
defparam \syif.store[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y73_N8
cycloneive_io_ibuf \syif.store[1]~input (
	.i(\syif.store [1]),
	.ibar(gnd),
	.o(\syif.store[1]~input_o ));
// synopsys translate_off
defparam \syif.store[1]~input .bus_hold = "false";
defparam \syif.store[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N15
cycloneive_io_ibuf \syif.store[2]~input (
	.i(\syif.store [2]),
	.ibar(gnd),
	.o(\syif.store[2]~input_o ));
// synopsys translate_off
defparam \syif.store[2]~input .bus_hold = "false";
defparam \syif.store[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N8
cycloneive_io_ibuf \syif.store[3]~input (
	.i(\syif.store [3]),
	.ibar(gnd),
	.o(\syif.store[3]~input_o ));
// synopsys translate_off
defparam \syif.store[3]~input .bus_hold = "false";
defparam \syif.store[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N8
cycloneive_io_ibuf \syif.store[4]~input (
	.i(\syif.store [4]),
	.ibar(gnd),
	.o(\syif.store[4]~input_o ));
// synopsys translate_off
defparam \syif.store[4]~input .bus_hold = "false";
defparam \syif.store[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N15
cycloneive_io_ibuf \syif.store[5]~input (
	.i(\syif.store [5]),
	.ibar(gnd),
	.o(\syif.store[5]~input_o ));
// synopsys translate_off
defparam \syif.store[5]~input .bus_hold = "false";
defparam \syif.store[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N1
cycloneive_io_ibuf \syif.store[6]~input (
	.i(\syif.store [6]),
	.ibar(gnd),
	.o(\syif.store[6]~input_o ));
// synopsys translate_off
defparam \syif.store[6]~input .bus_hold = "false";
defparam \syif.store[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N1
cycloneive_io_ibuf \syif.store[7]~input (
	.i(\syif.store [7]),
	.ibar(gnd),
	.o(\syif.store[7]~input_o ));
// synopsys translate_off
defparam \syif.store[7]~input .bus_hold = "false";
defparam \syif.store[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N15
cycloneive_io_ibuf \syif.store[8]~input (
	.i(\syif.store [8]),
	.ibar(gnd),
	.o(\syif.store[8]~input_o ));
// synopsys translate_off
defparam \syif.store[8]~input .bus_hold = "false";
defparam \syif.store[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y34_N15
cycloneive_io_ibuf \syif.store[9]~input (
	.i(\syif.store [9]),
	.ibar(gnd),
	.o(\syif.store[9]~input_o ));
// synopsys translate_off
defparam \syif.store[9]~input .bus_hold = "false";
defparam \syif.store[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N15
cycloneive_io_ibuf \syif.store[10]~input (
	.i(\syif.store [10]),
	.ibar(gnd),
	.o(\syif.store[10]~input_o ));
// synopsys translate_off
defparam \syif.store[10]~input .bus_hold = "false";
defparam \syif.store[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N8
cycloneive_io_ibuf \syif.store[11]~input (
	.i(\syif.store [11]),
	.ibar(gnd),
	.o(\syif.store[11]~input_o ));
// synopsys translate_off
defparam \syif.store[11]~input .bus_hold = "false";
defparam \syif.store[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X79_Y73_N1
cycloneive_io_ibuf \syif.store[12]~input (
	.i(\syif.store [12]),
	.ibar(gnd),
	.o(\syif.store[12]~input_o ));
// synopsys translate_off
defparam \syif.store[12]~input .bus_hold = "false";
defparam \syif.store[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N1
cycloneive_io_ibuf \syif.store[13]~input (
	.i(\syif.store [13]),
	.ibar(gnd),
	.o(\syif.store[13]~input_o ));
// synopsys translate_off
defparam \syif.store[13]~input .bus_hold = "false";
defparam \syif.store[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N8
cycloneive_io_ibuf \syif.store[14]~input (
	.i(\syif.store [14]),
	.ibar(gnd),
	.o(\syif.store[14]~input_o ));
// synopsys translate_off
defparam \syif.store[14]~input .bus_hold = "false";
defparam \syif.store[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y73_N22
cycloneive_io_ibuf \syif.store[15]~input (
	.i(\syif.store [15]),
	.ibar(gnd),
	.o(\syif.store[15]~input_o ));
// synopsys translate_off
defparam \syif.store[15]~input .bus_hold = "false";
defparam \syif.store[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y35_N22
cycloneive_io_ibuf \syif.store[16]~input (
	.i(\syif.store [16]),
	.ibar(gnd),
	.o(\syif.store[16]~input_o ));
// synopsys translate_off
defparam \syif.store[16]~input .bus_hold = "false";
defparam \syif.store[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N15
cycloneive_io_ibuf \syif.store[17]~input (
	.i(\syif.store [17]),
	.ibar(gnd),
	.o(\syif.store[17]~input_o ));
// synopsys translate_off
defparam \syif.store[17]~input .bus_hold = "false";
defparam \syif.store[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N8
cycloneive_io_ibuf \syif.store[18]~input (
	.i(\syif.store [18]),
	.ibar(gnd),
	.o(\syif.store[18]~input_o ));
// synopsys translate_off
defparam \syif.store[18]~input .bus_hold = "false";
defparam \syif.store[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y73_N1
cycloneive_io_ibuf \syif.store[19]~input (
	.i(\syif.store [19]),
	.ibar(gnd),
	.o(\syif.store[19]~input_o ));
// synopsys translate_off
defparam \syif.store[19]~input .bus_hold = "false";
defparam \syif.store[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N8
cycloneive_io_ibuf \syif.store[20]~input (
	.i(\syif.store [20]),
	.ibar(gnd),
	.o(\syif.store[20]~input_o ));
// synopsys translate_off
defparam \syif.store[20]~input .bus_hold = "false";
defparam \syif.store[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y34_N22
cycloneive_io_ibuf \syif.store[21]~input (
	.i(\syif.store [21]),
	.ibar(gnd),
	.o(\syif.store[21]~input_o ));
// synopsys translate_off
defparam \syif.store[21]~input .bus_hold = "false";
defparam \syif.store[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N1
cycloneive_io_ibuf \syif.store[22]~input (
	.i(\syif.store [22]),
	.ibar(gnd),
	.o(\syif.store[22]~input_o ));
// synopsys translate_off
defparam \syif.store[22]~input .bus_hold = "false";
defparam \syif.store[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N22
cycloneive_io_ibuf \syif.store[23]~input (
	.i(\syif.store [23]),
	.ibar(gnd),
	.o(\syif.store[23]~input_o ));
// synopsys translate_off
defparam \syif.store[23]~input .bus_hold = "false";
defparam \syif.store[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N15
cycloneive_io_ibuf \syif.store[24]~input (
	.i(\syif.store [24]),
	.ibar(gnd),
	.o(\syif.store[24]~input_o ));
// synopsys translate_off
defparam \syif.store[24]~input .bus_hold = "false";
defparam \syif.store[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y73_N15
cycloneive_io_ibuf \syif.store[25]~input (
	.i(\syif.store [25]),
	.ibar(gnd),
	.o(\syif.store[25]~input_o ));
// synopsys translate_off
defparam \syif.store[25]~input .bus_hold = "false";
defparam \syif.store[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N1
cycloneive_io_ibuf \syif.store[26]~input (
	.i(\syif.store [26]),
	.ibar(gnd),
	.o(\syif.store[26]~input_o ));
// synopsys translate_off
defparam \syif.store[26]~input .bus_hold = "false";
defparam \syif.store[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y33_N1
cycloneive_io_ibuf \syif.store[27]~input (
	.i(\syif.store [27]),
	.ibar(gnd),
	.o(\syif.store[27]~input_o ));
// synopsys translate_off
defparam \syif.store[27]~input .bus_hold = "false";
defparam \syif.store[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X79_Y73_N8
cycloneive_io_ibuf \syif.store[28]~input (
	.i(\syif.store [28]),
	.ibar(gnd),
	.o(\syif.store[28]~input_o ));
// synopsys translate_off
defparam \syif.store[28]~input .bus_hold = "false";
defparam \syif.store[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N1
cycloneive_io_ibuf \syif.store[29]~input (
	.i(\syif.store [29]),
	.ibar(gnd),
	.o(\syif.store[29]~input_o ));
// synopsys translate_off
defparam \syif.store[29]~input .bus_hold = "false";
defparam \syif.store[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N8
cycloneive_io_ibuf \syif.store[30]~input (
	.i(\syif.store [30]),
	.ibar(gnd),
	.o(\syif.store[30]~input_o ));
// synopsys translate_off
defparam \syif.store[30]~input .bus_hold = "false";
defparam \syif.store[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N22
cycloneive_io_ibuf \syif.store[31]~input (
	.i(\syif.store [31]),
	.ibar(gnd),
	.o(\syif.store[31]~input_o ));
// synopsys translate_off
defparam \syif.store[31]~input .bus_hold = "false";
defparam \syif.store[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: CLKCTRL_G4
cycloneive_clkctrl \altera_internal_jtag~TCKUTAPclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\altera_internal_jtag~TCKUTAP }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ));
// synopsys translate_off
defparam \altera_internal_jtag~TCKUTAPclkctrl .clock_type = "global clock";
defparam \altera_internal_jtag~TCKUTAPclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G10
cycloneive_clkctrl \CPUCLK~clkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CPUCLK~q }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CPUCLK~clkctrl_outclk ));
// synopsys translate_off
defparam \CPUCLK~clkctrl .clock_type = "global clock";
defparam \CPUCLK~clkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G1
cycloneive_clkctrl \nRST~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\nRST~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\nRST~inputclkctrl_outclk ));
// synopsys translate_off
defparam \nRST~inputclkctrl .clock_type = "global clock";
defparam \nRST~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G2
cycloneive_clkctrl \CLK~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CLK~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CLK~inputclkctrl_outclk ));
// synopsys translate_off
defparam \CLK~inputclkctrl .clock_type = "global clock";
defparam \CLK~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: LCCOMB_X45_Y41_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y41_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y41_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N23
cycloneive_io_obuf \syif.halt~output (
	.i(\CPU|DP|dpif.halt~q ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.halt ),
	.obar());
// synopsys translate_off
defparam \syif.halt~output .bus_hold = "false";
defparam \syif.halt~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N9
cycloneive_io_obuf \syif.load[0]~output (
	.i(\RAM|ramif.ramload[0]~0_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [0]),
	.obar());
// synopsys translate_off
defparam \syif.load[0]~output .bus_hold = "false";
defparam \syif.load[0]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y42_N2
cycloneive_io_obuf \syif.load[1]~output (
	.i(\RAM|ramif.ramload[1]~1_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [1]),
	.obar());
// synopsys translate_off
defparam \syif.load[1]~output .bus_hold = "false";
defparam \syif.load[1]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N23
cycloneive_io_obuf \syif.load[2]~output (
	.i(\RAM|ramif.ramload[2]~2_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [2]),
	.obar());
// synopsys translate_off
defparam \syif.load[2]~output .bus_hold = "false";
defparam \syif.load[2]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y41_N9
cycloneive_io_obuf \syif.load[3]~output (
	.i(\RAM|ramif.ramload[3]~3_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [3]),
	.obar());
// synopsys translate_off
defparam \syif.load[3]~output .bus_hold = "false";
defparam \syif.load[3]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y0_N23
cycloneive_io_obuf \syif.load[4]~output (
	.i(\RAM|ramif.ramload[4]~4_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [4]),
	.obar());
// synopsys translate_off
defparam \syif.load[4]~output .bus_hold = "false";
defparam \syif.load[4]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N23
cycloneive_io_obuf \syif.load[5]~output (
	.i(\RAM|ramif.ramload[5]~5_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [5]),
	.obar());
// synopsys translate_off
defparam \syif.load[5]~output .bus_hold = "false";
defparam \syif.load[5]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X83_Y73_N2
cycloneive_io_obuf \syif.load[6]~output (
	.i(\RAM|ramif.ramload[6]~6_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [6]),
	.obar());
// synopsys translate_off
defparam \syif.load[6]~output .bus_hold = "false";
defparam \syif.load[6]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X72_Y73_N16
cycloneive_io_obuf \syif.load[7]~output (
	.i(\RAM|ramif.ramload[7]~7_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [7]),
	.obar());
// synopsys translate_off
defparam \syif.load[7]~output .bus_hold = "false";
defparam \syif.load[7]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X74_Y73_N23
cycloneive_io_obuf \syif.load[8]~output (
	.i(\RAM|ramif.ramload[8]~8_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [8]),
	.obar());
// synopsys translate_off
defparam \syif.load[8]~output .bus_hold = "false";
defparam \syif.load[8]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X74_Y0_N23
cycloneive_io_obuf \syif.load[9]~output (
	.i(\RAM|ramif.ramload[9]~9_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [9]),
	.obar());
// synopsys translate_off
defparam \syif.load[9]~output .bus_hold = "false";
defparam \syif.load[9]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y40_N9
cycloneive_io_obuf \syif.load[10]~output (
	.i(\RAM|ramif.ramload[10]~10_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [10]),
	.obar());
// synopsys translate_off
defparam \syif.load[10]~output .bus_hold = "false";
defparam \syif.load[10]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y73_N23
cycloneive_io_obuf \syif.load[11]~output (
	.i(\RAM|ramif.ramload[11]~11_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [11]),
	.obar());
// synopsys translate_off
defparam \syif.load[11]~output .bus_hold = "false";
defparam \syif.load[11]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X81_Y73_N2
cycloneive_io_obuf \syif.load[12]~output (
	.i(\RAM|ramif.ramload[12]~12_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [12]),
	.obar());
// synopsys translate_off
defparam \syif.load[12]~output .bus_hold = "false";
defparam \syif.load[12]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X81_Y73_N16
cycloneive_io_obuf \syif.load[13]~output (
	.i(\RAM|ramif.ramload[13]~13_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [13]),
	.obar());
// synopsys translate_off
defparam \syif.load[13]~output .bus_hold = "false";
defparam \syif.load[13]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y73_N16
cycloneive_io_obuf \syif.load[14]~output (
	.i(\RAM|ramif.ramload[14]~14_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [14]),
	.obar());
// synopsys translate_off
defparam \syif.load[14]~output .bus_hold = "false";
defparam \syif.load[14]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N16
cycloneive_io_obuf \syif.load[15]~output (
	.i(\RAM|ramif.ramload[15]~15_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [15]),
	.obar());
// synopsys translate_off
defparam \syif.load[15]~output .bus_hold = "false";
defparam \syif.load[15]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y73_N9
cycloneive_io_obuf \syif.load[16]~output (
	.i(\RAM|ramif.ramload[16]~16_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [16]),
	.obar());
// synopsys translate_off
defparam \syif.load[16]~output .bus_hold = "false";
defparam \syif.load[16]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N2
cycloneive_io_obuf \syif.load[17]~output (
	.i(\RAM|ramif.ramload[17]~17_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [17]),
	.obar());
// synopsys translate_off
defparam \syif.load[17]~output .bus_hold = "false";
defparam \syif.load[17]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y73_N2
cycloneive_io_obuf \syif.load[18]~output (
	.i(\RAM|ramif.ramload[18]~18_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [18]),
	.obar());
// synopsys translate_off
defparam \syif.load[18]~output .bus_hold = "false";
defparam \syif.load[18]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y0_N16
cycloneive_io_obuf \syif.load[19]~output (
	.i(\RAM|ramif.ramload[19]~19_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [19]),
	.obar());
// synopsys translate_off
defparam \syif.load[19]~output .bus_hold = "false";
defparam \syif.load[19]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N16
cycloneive_io_obuf \syif.load[20]~output (
	.i(\RAM|ramif.ramload[20]~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [20]),
	.obar());
// synopsys translate_off
defparam \syif.load[20]~output .bus_hold = "false";
defparam \syif.load[20]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N16
cycloneive_io_obuf \syif.load[21]~output (
	.i(\RAM|ramif.ramload[21]~21_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [21]),
	.obar());
// synopsys translate_off
defparam \syif.load[21]~output .bus_hold = "false";
defparam \syif.load[21]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y0_N9
cycloneive_io_obuf \syif.load[22]~output (
	.i(\RAM|ramif.ramload[22]~22_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [22]),
	.obar());
// synopsys translate_off
defparam \syif.load[22]~output .bus_hold = "false";
defparam \syif.load[22]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y73_N16
cycloneive_io_obuf \syif.load[23]~output (
	.i(\RAM|ramif.ramload[23]~23_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [23]),
	.obar());
// synopsys translate_off
defparam \syif.load[23]~output .bus_hold = "false";
defparam \syif.load[23]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y0_N2
cycloneive_io_obuf \syif.load[24]~output (
	.i(\RAM|ramif.ramload[24]~24_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [24]),
	.obar());
// synopsys translate_off
defparam \syif.load[24]~output .bus_hold = "false";
defparam \syif.load[24]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y73_N2
cycloneive_io_obuf \syif.load[25]~output (
	.i(\RAM|ramif.ramload[25]~25_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [25]),
	.obar());
// synopsys translate_off
defparam \syif.load[25]~output .bus_hold = "false";
defparam \syif.load[25]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N9
cycloneive_io_obuf \syif.load[26]~output (
	.i(\RAM|ramif.ramload[26]~26_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [26]),
	.obar());
// synopsys translate_off
defparam \syif.load[26]~output .bus_hold = "false";
defparam \syif.load[26]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N2
cycloneive_io_obuf \syif.load[27]~output (
	.i(\RAM|ramif.ramload[27]~27_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [27]),
	.obar());
// synopsys translate_off
defparam \syif.load[27]~output .bus_hold = "false";
defparam \syif.load[27]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X81_Y73_N23
cycloneive_io_obuf \syif.load[28]~output (
	.i(\RAM|ramif.ramload[28]~28_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [28]),
	.obar());
// synopsys translate_off
defparam \syif.load[28]~output .bus_hold = "false";
defparam \syif.load[28]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N23
cycloneive_io_obuf \syif.load[29]~output (
	.i(\RAM|ramif.ramload[29]~29_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [29]),
	.obar());
// synopsys translate_off
defparam \syif.load[29]~output .bus_hold = "false";
defparam \syif.load[29]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N16
cycloneive_io_obuf \syif.load[30]~output (
	.i(\RAM|ramif.ramload[30]~30_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [30]),
	.obar());
// synopsys translate_off
defparam \syif.load[30]~output .bus_hold = "false";
defparam \syif.load[30]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N2
cycloneive_io_obuf \syif.load[31]~output (
	.i(\RAM|ramif.ramload[31]~31_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [31]),
	.obar());
// synopsys translate_off
defparam \syif.load[31]~output .bus_hold = "false";
defparam \syif.load[31]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y37_N1
cycloneive_io_obuf \altera_reserved_tdo~output (
	.i(\altera_internal_jtag~TDO ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(altera_reserved_tdo),
	.obar());
// synopsys translate_off
defparam \altera_reserved_tdo~output .bus_hold = "false";
defparam \altera_reserved_tdo~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOIBUF_X0_Y38_N1
cycloneive_io_ibuf \altera_reserved_tms~input (
	.i(altera_reserved_tms),
	.ibar(gnd),
	.o(\altera_reserved_tms~input_o ));
// synopsys translate_off
defparam \altera_reserved_tms~input .bus_hold = "false";
defparam \altera_reserved_tms~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y39_N1
cycloneive_io_ibuf \altera_reserved_tck~input (
	.i(altera_reserved_tck),
	.ibar(gnd),
	.o(\altera_reserved_tck~input_o ));
// synopsys translate_off
defparam \altera_reserved_tck~input .bus_hold = "false";
defparam \altera_reserved_tck~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y40_N1
cycloneive_io_ibuf \altera_reserved_tdi~input (
	.i(altera_reserved_tdi),
	.ibar(gnd),
	.o(\altera_reserved_tdi~input_o ));
// synopsys translate_off
defparam \altera_reserved_tdi~input .bus_hold = "false";
defparam \altera_reserved_tdi~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h33CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y40_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .lut_mask = 16'h5500;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .lut_mask = 16'hFFFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .lut_mask = 16'hAA88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .lut_mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hAA88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .lut_mask = 16'hAA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .lut_mask = 16'hEE00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .lut_mask = 16'hFFFD;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .lut_mask = 16'hAAA8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y40_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .lut_mask = 16'h0C0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y40_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .lut_mask = 16'h5AF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y40_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .lut_mask = 16'h5575;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y40_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y39_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y39_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .lut_mask = 16'h0010;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .lut_mask = 16'h0800;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .lut_mask = 16'hFFFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y42_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .lut_mask = 16'hAAEA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y42_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .lut_mask = 16'h0200;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y39_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .lut_mask = 16'hC30C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .lut_mask = 16'hC3C3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X45_Y42_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .lut_mask = 16'hB3A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y42_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y42_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y42_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .lut_mask = 16'h1110;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .lut_mask = 16'h3320;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y40_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .lut_mask = 16'hFAF8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y42_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .lut_mask = 16'h0002;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .lut_mask = 16'hFF20;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y42_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .lut_mask = 16'hF022;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .lut_mask = 16'h4C4C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y42_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y42_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .lut_mask = 16'hAEAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y42_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .lut_mask = 16'h00F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .lut_mask = 16'hFCFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y41_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .lut_mask = 16'hFFCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y41_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .lut_mask = 16'h3300;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y41_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .lut_mask = 16'hFFCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y41_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y42_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .lut_mask = 16'hAAF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y42_N22
cycloneive_lcell_comb \~QIC_CREATED_GND~I (
// Equation(s):
// \~QIC_CREATED_GND~I_combout  = GND

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.cout());
// synopsys translate_off
defparam \~QIC_CREATED_GND~I .lut_mask = 16'h0000;
defparam \~QIC_CREATED_GND~I .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .lut_mask = 16'hAA88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .lut_mask = 16'h8880;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y41_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y41_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .lut_mask = 16'h50C2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .lut_mask = 16'hB4F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y41_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .lut_mask = 16'h0800;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .lut_mask = 16'h7430;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y41_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y40_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .lut_mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y40_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y42_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.asdata(\~QIC_CREATED_GND~I_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .lut_mask = 16'hFA50;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .lut_mask = 16'h0088;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .lut_mask = 16'h7430;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y41_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 (
	.dataa(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .lut_mask = 16'hBB88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y41_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 (
	.dataa(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .lut_mask = 16'hAFA0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y41_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .lut_mask = 16'hA808;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y41_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y41_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .lut_mask = 16'hCFC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y41_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y41_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 (
	.dataa(gnd),
	.datab(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .lut_mask = 16'hCFC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y41_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y41_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 (
	.dataa(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .lut_mask = 16'hAFA0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y41_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y41_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .lut_mask = 16'hFA50;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y41_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .lut_mask = 16'hAAE4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y41_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .lut_mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y41_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .lut_mask = 16'hAAE4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 .lut_mask = 16'hA505;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 .lut_mask = 16'h3CCF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y40_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .lut_mask = 16'hECA0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y40_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 .lut_mask = 16'h0003;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .lut_mask = 16'hFF10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y40_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X41_Y40_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .lut_mask = 16'h3C3C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X41_Y40_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5 .lut_mask = 16'h8000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y40_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .lut_mask = 16'h0080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .lut_mask = 16'h00C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y40_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y40_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y40_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y40_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y40_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y40_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y40_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .lut_mask = 16'h0020;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y40_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y40_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7 .lut_mask = 16'h0002;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y40_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .lut_mask = 16'hEFC8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y40_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y40_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 .lut_mask = 16'hF0CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y40_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .lut_mask = 16'hDD88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y40_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y40_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y40_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y40_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y40_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y40_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y40_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .lut_mask = 16'h33FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y40_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .lut_mask = 16'hFC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y40_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y40_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y40_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y40_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y41_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .lut_mask = 16'h15BB;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y41_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo (
	.clk(!\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X28_Y38_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X5_Y14_N0
cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y39_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline (
	dpifhalt,
	temp_aluResult_1,
	pccount_1,
	temp_dmemWEN,
	temp_dmemREN,
	temp_aluResult_0,
	pccount_0,
	temp_aluResult_2,
	pccount_2,
	temp_aluResult_3,
	pccount_3,
	temp_aluResult_5,
	pccount_5,
	temp_aluResult_4,
	pccount_4,
	temp_aluResult_7,
	pccount_7,
	temp_aluResult_6,
	pccount_6,
	temp_aluResult_9,
	pccount_9,
	temp_aluResult_8,
	pccount_8,
	temp_aluResult_11,
	pccount_11,
	temp_aluResult_10,
	pccount_10,
	temp_aluResult_13,
	pccount_13,
	temp_aluResult_12,
	pccount_12,
	temp_aluResult_15,
	pccount_15,
	temp_aluResult_14,
	pccount_14,
	temp_aluResult_17,
	pccount_17,
	temp_aluResult_16,
	pccount_16,
	temp_aluResult_19,
	pccount_19,
	temp_aluResult_18,
	pccount_18,
	temp_aluResult_20,
	pccount_20,
	temp_aluResult_21,
	pccount_21,
	temp_aluResult_23,
	pccount_23,
	temp_aluResult_22,
	pccount_22,
	temp_aluResult_25,
	pccount_25,
	temp_aluResult_24,
	pccount_24,
	temp_aluResult_26,
	pccount_26,
	temp_aluResult_27,
	pccount_27,
	temp_aluResult_29,
	pccount_29,
	temp_aluResult_28,
	pccount_28,
	temp_aluResult_31,
	pccount_31,
	temp_aluResult_30,
	pccount_30,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	temp_rdat2_0,
	temp_rdat2_1,
	temp_rdat2_2,
	temp_rdat2_3,
	temp_rdat2_4,
	temp_rdat2_5,
	temp_rdat2_6,
	temp_rdat2_7,
	temp_rdat2_8,
	temp_rdat2_9,
	temp_rdat2_10,
	temp_rdat2_11,
	temp_rdat2_12,
	temp_rdat2_13,
	temp_rdat2_14,
	temp_rdat2_15,
	temp_rdat2_16,
	temp_rdat2_17,
	temp_rdat2_18,
	temp_rdat2_19,
	temp_rdat2_20,
	temp_rdat2_21,
	temp_rdat2_22,
	temp_rdat2_23,
	temp_rdat2_24,
	temp_rdat2_25,
	temp_rdat2_26,
	temp_rdat2_27,
	temp_rdat2_28,
	temp_rdat2_29,
	temp_rdat2_30,
	temp_rdat2_31,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	dpifhalt;
output 	temp_aluResult_1;
output 	pccount_1;
output 	temp_dmemWEN;
output 	temp_dmemREN;
output 	temp_aluResult_0;
output 	pccount_0;
output 	temp_aluResult_2;
output 	pccount_2;
output 	temp_aluResult_3;
output 	pccount_3;
output 	temp_aluResult_5;
output 	pccount_5;
output 	temp_aluResult_4;
output 	pccount_4;
output 	temp_aluResult_7;
output 	pccount_7;
output 	temp_aluResult_6;
output 	pccount_6;
output 	temp_aluResult_9;
output 	pccount_9;
output 	temp_aluResult_8;
output 	pccount_8;
output 	temp_aluResult_11;
output 	pccount_11;
output 	temp_aluResult_10;
output 	pccount_10;
output 	temp_aluResult_13;
output 	pccount_13;
output 	temp_aluResult_12;
output 	pccount_12;
output 	temp_aluResult_15;
output 	pccount_15;
output 	temp_aluResult_14;
output 	pccount_14;
output 	temp_aluResult_17;
output 	pccount_17;
output 	temp_aluResult_16;
output 	pccount_16;
output 	temp_aluResult_19;
output 	pccount_19;
output 	temp_aluResult_18;
output 	pccount_18;
output 	temp_aluResult_20;
output 	pccount_20;
output 	temp_aluResult_21;
output 	pccount_21;
output 	temp_aluResult_23;
output 	pccount_23;
output 	temp_aluResult_22;
output 	pccount_22;
output 	temp_aluResult_25;
output 	pccount_25;
output 	temp_aluResult_24;
output 	pccount_24;
output 	temp_aluResult_26;
output 	pccount_26;
output 	temp_aluResult_27;
output 	pccount_27;
output 	temp_aluResult_29;
output 	pccount_29;
output 	temp_aluResult_28;
output 	pccount_28;
output 	temp_aluResult_31;
output 	pccount_31;
output 	temp_aluResult_30;
output 	pccount_30;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	temp_rdat2_0;
output 	temp_rdat2_1;
output 	temp_rdat2_2;
output 	temp_rdat2_3;
output 	temp_rdat2_4;
output 	temp_rdat2_5;
output 	temp_rdat2_6;
output 	temp_rdat2_7;
output 	temp_rdat2_8;
output 	temp_rdat2_9;
output 	temp_rdat2_10;
output 	temp_rdat2_11;
output 	temp_rdat2_12;
output 	temp_rdat2_13;
output 	temp_rdat2_14;
output 	temp_rdat2_15;
output 	temp_rdat2_16;
output 	temp_rdat2_17;
output 	temp_rdat2_18;
output 	temp_rdat2_19;
output 	temp_rdat2_20;
output 	temp_rdat2_21;
output 	temp_rdat2_22;
output 	temp_rdat2_23;
output 	temp_rdat2_24;
output 	temp_rdat2_25;
output 	temp_rdat2_26;
output 	temp_rdat2_27;
output 	temp_rdat2_28;
output 	temp_rdat2_29;
output 	temp_rdat2_30;
output 	temp_rdat2_31;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \CC|ccif.iwait[0]~0_combout ;


memory_control CC(
	.temp_dmemWEN(temp_dmemWEN),
	.temp_dmemREN(temp_dmemREN),
	.always1(always1),
	.ccifiwait_0(\CC|ccif.iwait[0]~0_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

datapath DP(
	.dpifhalt(dpifhalt),
	.temp_aluResult_1(temp_aluResult_1),
	.pccount_1(pccount_1),
	.temp_dmemWEN(temp_dmemWEN),
	.temp_dmemREN(temp_dmemREN),
	.temp_aluResult_0(temp_aluResult_0),
	.pccount_0(pccount_0),
	.temp_aluResult_2(temp_aluResult_2),
	.pccount_2(pccount_2),
	.temp_aluResult_3(temp_aluResult_3),
	.pccount_3(pccount_3),
	.temp_aluResult_5(temp_aluResult_5),
	.pccount_5(pccount_5),
	.temp_aluResult_4(temp_aluResult_4),
	.pccount_4(pccount_4),
	.temp_aluResult_7(temp_aluResult_7),
	.pccount_7(pccount_7),
	.temp_aluResult_6(temp_aluResult_6),
	.pccount_6(pccount_6),
	.temp_aluResult_9(temp_aluResult_9),
	.pccount_9(pccount_9),
	.temp_aluResult_8(temp_aluResult_8),
	.pccount_8(pccount_8),
	.temp_aluResult_11(temp_aluResult_11),
	.pccount_11(pccount_11),
	.temp_aluResult_10(temp_aluResult_10),
	.pccount_10(pccount_10),
	.temp_aluResult_13(temp_aluResult_13),
	.pccount_13(pccount_13),
	.temp_aluResult_12(temp_aluResult_12),
	.pccount_12(pccount_12),
	.temp_aluResult_15(temp_aluResult_15),
	.pccount_15(pccount_15),
	.temp_aluResult_14(temp_aluResult_14),
	.pccount_14(pccount_14),
	.temp_aluResult_17(temp_aluResult_17),
	.pccount_17(pccount_17),
	.temp_aluResult_16(temp_aluResult_16),
	.pccount_16(pccount_16),
	.temp_aluResult_19(temp_aluResult_19),
	.pccount_19(pccount_19),
	.temp_aluResult_18(temp_aluResult_18),
	.pccount_18(pccount_18),
	.temp_aluResult_20(temp_aluResult_20),
	.pccount_20(pccount_20),
	.temp_aluResult_21(temp_aluResult_21),
	.pccount_21(pccount_21),
	.temp_aluResult_23(temp_aluResult_23),
	.pccount_23(pccount_23),
	.temp_aluResult_22(temp_aluResult_22),
	.pccount_22(pccount_22),
	.temp_aluResult_25(temp_aluResult_25),
	.pccount_25(pccount_25),
	.temp_aluResult_24(temp_aluResult_24),
	.pccount_24(pccount_24),
	.temp_aluResult_26(temp_aluResult_26),
	.pccount_26(pccount_26),
	.temp_aluResult_27(temp_aluResult_27),
	.pccount_27(pccount_27),
	.temp_aluResult_29(temp_aluResult_29),
	.pccount_29(pccount_29),
	.temp_aluResult_28(temp_aluResult_28),
	.pccount_28(pccount_28),
	.temp_aluResult_31(temp_aluResult_31),
	.pccount_31(pccount_31),
	.temp_aluResult_30(temp_aluResult_30),
	.pccount_30(pccount_30),
	.always1(always1),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.temp_rdat2_0(temp_rdat2_0),
	.ccifiwait_0(\CC|ccif.iwait[0]~0_combout ),
	.temp_rdat2_1(temp_rdat2_1),
	.temp_rdat2_2(temp_rdat2_2),
	.temp_rdat2_3(temp_rdat2_3),
	.temp_rdat2_4(temp_rdat2_4),
	.temp_rdat2_5(temp_rdat2_5),
	.temp_rdat2_6(temp_rdat2_6),
	.temp_rdat2_7(temp_rdat2_7),
	.temp_rdat2_8(temp_rdat2_8),
	.temp_rdat2_9(temp_rdat2_9),
	.temp_rdat2_10(temp_rdat2_10),
	.temp_rdat2_11(temp_rdat2_11),
	.temp_rdat2_12(temp_rdat2_12),
	.temp_rdat2_13(temp_rdat2_13),
	.temp_rdat2_14(temp_rdat2_14),
	.temp_rdat2_15(temp_rdat2_15),
	.temp_rdat2_16(temp_rdat2_16),
	.temp_rdat2_17(temp_rdat2_17),
	.temp_rdat2_18(temp_rdat2_18),
	.temp_rdat2_19(temp_rdat2_19),
	.temp_rdat2_20(temp_rdat2_20),
	.temp_rdat2_21(temp_rdat2_21),
	.temp_rdat2_22(temp_rdat2_22),
	.temp_rdat2_23(temp_rdat2_23),
	.temp_rdat2_24(temp_rdat2_24),
	.temp_rdat2_25(temp_rdat2_25),
	.temp_rdat2_26(temp_rdat2_26),
	.temp_rdat2_27(temp_rdat2_27),
	.temp_rdat2_28(temp_rdat2_28),
	.temp_rdat2_29(temp_rdat2_29),
	.temp_rdat2_30(temp_rdat2_30),
	.temp_rdat2_31(temp_rdat2_31),
	.CPUCLK(CPUCLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module datapath (
	dpifhalt,
	temp_aluResult_1,
	pccount_1,
	temp_dmemWEN,
	temp_dmemREN,
	temp_aluResult_0,
	pccount_0,
	temp_aluResult_2,
	pccount_2,
	temp_aluResult_3,
	pccount_3,
	temp_aluResult_5,
	pccount_5,
	temp_aluResult_4,
	pccount_4,
	temp_aluResult_7,
	pccount_7,
	temp_aluResult_6,
	pccount_6,
	temp_aluResult_9,
	pccount_9,
	temp_aluResult_8,
	pccount_8,
	temp_aluResult_11,
	pccount_11,
	temp_aluResult_10,
	pccount_10,
	temp_aluResult_13,
	pccount_13,
	temp_aluResult_12,
	pccount_12,
	temp_aluResult_15,
	pccount_15,
	temp_aluResult_14,
	pccount_14,
	temp_aluResult_17,
	pccount_17,
	temp_aluResult_16,
	pccount_16,
	temp_aluResult_19,
	pccount_19,
	temp_aluResult_18,
	pccount_18,
	temp_aluResult_20,
	pccount_20,
	temp_aluResult_21,
	pccount_21,
	temp_aluResult_23,
	pccount_23,
	temp_aluResult_22,
	pccount_22,
	temp_aluResult_25,
	pccount_25,
	temp_aluResult_24,
	pccount_24,
	temp_aluResult_26,
	pccount_26,
	temp_aluResult_27,
	pccount_27,
	temp_aluResult_29,
	pccount_29,
	temp_aluResult_28,
	pccount_28,
	temp_aluResult_31,
	pccount_31,
	temp_aluResult_30,
	pccount_30,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	temp_rdat2_0,
	ccifiwait_0,
	temp_rdat2_1,
	temp_rdat2_2,
	temp_rdat2_3,
	temp_rdat2_4,
	temp_rdat2_5,
	temp_rdat2_6,
	temp_rdat2_7,
	temp_rdat2_8,
	temp_rdat2_9,
	temp_rdat2_10,
	temp_rdat2_11,
	temp_rdat2_12,
	temp_rdat2_13,
	temp_rdat2_14,
	temp_rdat2_15,
	temp_rdat2_16,
	temp_rdat2_17,
	temp_rdat2_18,
	temp_rdat2_19,
	temp_rdat2_20,
	temp_rdat2_21,
	temp_rdat2_22,
	temp_rdat2_23,
	temp_rdat2_24,
	temp_rdat2_25,
	temp_rdat2_26,
	temp_rdat2_27,
	temp_rdat2_28,
	temp_rdat2_29,
	temp_rdat2_30,
	temp_rdat2_31,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	dpifhalt;
output 	temp_aluResult_1;
output 	pccount_1;
output 	temp_dmemWEN;
output 	temp_dmemREN;
output 	temp_aluResult_0;
output 	pccount_0;
output 	temp_aluResult_2;
output 	pccount_2;
output 	temp_aluResult_3;
output 	pccount_3;
output 	temp_aluResult_5;
output 	pccount_5;
output 	temp_aluResult_4;
output 	pccount_4;
output 	temp_aluResult_7;
output 	pccount_7;
output 	temp_aluResult_6;
output 	pccount_6;
output 	temp_aluResult_9;
output 	pccount_9;
output 	temp_aluResult_8;
output 	pccount_8;
output 	temp_aluResult_11;
output 	pccount_11;
output 	temp_aluResult_10;
output 	pccount_10;
output 	temp_aluResult_13;
output 	pccount_13;
output 	temp_aluResult_12;
output 	pccount_12;
output 	temp_aluResult_15;
output 	pccount_15;
output 	temp_aluResult_14;
output 	pccount_14;
output 	temp_aluResult_17;
output 	pccount_17;
output 	temp_aluResult_16;
output 	pccount_16;
output 	temp_aluResult_19;
output 	pccount_19;
output 	temp_aluResult_18;
output 	pccount_18;
output 	temp_aluResult_20;
output 	pccount_20;
output 	temp_aluResult_21;
output 	pccount_21;
output 	temp_aluResult_23;
output 	pccount_23;
output 	temp_aluResult_22;
output 	pccount_22;
output 	temp_aluResult_25;
output 	pccount_25;
output 	temp_aluResult_24;
output 	pccount_24;
output 	temp_aluResult_26;
output 	pccount_26;
output 	temp_aluResult_27;
output 	pccount_27;
output 	temp_aluResult_29;
output 	pccount_29;
output 	temp_aluResult_28;
output 	pccount_28;
output 	temp_aluResult_31;
output 	pccount_31;
output 	temp_aluResult_30;
output 	pccount_30;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	temp_rdat2_0;
input 	ccifiwait_0;
output 	temp_rdat2_1;
output 	temp_rdat2_2;
output 	temp_rdat2_3;
output 	temp_rdat2_4;
output 	temp_rdat2_5;
output 	temp_rdat2_6;
output 	temp_rdat2_7;
output 	temp_rdat2_8;
output 	temp_rdat2_9;
output 	temp_rdat2_10;
output 	temp_rdat2_11;
output 	temp_rdat2_12;
output 	temp_rdat2_13;
output 	temp_rdat2_14;
output 	temp_rdat2_15;
output 	temp_rdat2_16;
output 	temp_rdat2_17;
output 	temp_rdat2_18;
output 	temp_rdat2_19;
output 	temp_rdat2_20;
output 	temp_rdat2_21;
output 	temp_rdat2_22;
output 	temp_rdat2_23;
output 	temp_rdat2_24;
output 	temp_rdat2_25;
output 	temp_rdat2_26;
output 	temp_rdat2_27;
output 	temp_rdat2_28;
output 	temp_rdat2_29;
output 	temp_rdat2_30;
output 	temp_rdat2_31;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \EXMEM|temp_zeroFlag~q ;
wire \branch_count_output[2]~1 ;
wire \branch_count_output[2]~0_combout ;
wire \pc_count_four_output[2]~1 ;
wire \pc_count_four_output[2]~0_combout ;
wire \pc_count_four_output[3]~3 ;
wire \pc_count_four_output[3]~2_combout ;
wire \branch_count_output[3]~3 ;
wire \branch_count_output[3]~2_combout ;
wire \pc_count_four_output[4]~5 ;
wire \pc_count_four_output[4]~4_combout ;
wire \pc_count_four_output[5]~7 ;
wire \pc_count_four_output[5]~6_combout ;
wire \branch_count_output[4]~5 ;
wire \branch_count_output[4]~4_combout ;
wire \branch_count_output[5]~7 ;
wire \branch_count_output[5]~6_combout ;
wire \pc_count_four_output[6]~9 ;
wire \pc_count_four_output[6]~8_combout ;
wire \pc_count_four_output[7]~11 ;
wire \pc_count_four_output[7]~10_combout ;
wire \branch_count_output[6]~9 ;
wire \branch_count_output[6]~8_combout ;
wire \branch_count_output[7]~11 ;
wire \branch_count_output[7]~10_combout ;
wire \pc_count_four_output[8]~13 ;
wire \pc_count_four_output[8]~12_combout ;
wire \pc_count_four_output[9]~15 ;
wire \pc_count_four_output[9]~14_combout ;
wire \branch_count_output[8]~13 ;
wire \branch_count_output[8]~12_combout ;
wire \branch_count_output[9]~15 ;
wire \branch_count_output[9]~14_combout ;
wire \pc_count_four_output[10]~17 ;
wire \pc_count_four_output[10]~16_combout ;
wire \pc_count_four_output[11]~19 ;
wire \pc_count_four_output[11]~18_combout ;
wire \branch_count_output[10]~17 ;
wire \branch_count_output[10]~16_combout ;
wire \branch_count_output[11]~19 ;
wire \branch_count_output[11]~18_combout ;
wire \pc_count_four_output[12]~21 ;
wire \pc_count_four_output[12]~20_combout ;
wire \pc_count_four_output[13]~23 ;
wire \pc_count_four_output[13]~22_combout ;
wire \branch_count_output[12]~21 ;
wire \branch_count_output[12]~20_combout ;
wire \branch_count_output[13]~23 ;
wire \branch_count_output[13]~22_combout ;
wire \pc_count_four_output[14]~25 ;
wire \pc_count_four_output[14]~24_combout ;
wire \pc_count_four_output[15]~27 ;
wire \pc_count_four_output[15]~26_combout ;
wire \branch_count_output[14]~25 ;
wire \branch_count_output[14]~24_combout ;
wire \branch_count_output[15]~27 ;
wire \branch_count_output[15]~26_combout ;
wire \pc_count_four_output[16]~29 ;
wire \pc_count_four_output[16]~28_combout ;
wire \pc_count_four_output[17]~31 ;
wire \pc_count_four_output[17]~30_combout ;
wire \branch_count_output[16]~29 ;
wire \branch_count_output[16]~28_combout ;
wire \branch_count_output[17]~31 ;
wire \branch_count_output[17]~30_combout ;
wire \pc_count_four_output[18]~33 ;
wire \pc_count_four_output[18]~32_combout ;
wire \pc_count_four_output[19]~35 ;
wire \pc_count_four_output[19]~34_combout ;
wire \branch_count_output[18]~33 ;
wire \branch_count_output[18]~32_combout ;
wire \branch_count_output[19]~35 ;
wire \branch_count_output[19]~34_combout ;
wire \branch_count_output[20]~37 ;
wire \branch_count_output[20]~36_combout ;
wire \pc_count_four_output[20]~37 ;
wire \pc_count_four_output[20]~36_combout ;
wire \pc_count_four_output[21]~39 ;
wire \pc_count_four_output[21]~38_combout ;
wire \branch_count_output[21]~39 ;
wire \branch_count_output[21]~38_combout ;
wire \pc_count_four_output[22]~41 ;
wire \pc_count_four_output[22]~40_combout ;
wire \pc_count_four_output[23]~43 ;
wire \pc_count_four_output[23]~42_combout ;
wire \branch_count_output[22]~41 ;
wire \branch_count_output[22]~40_combout ;
wire \branch_count_output[23]~43 ;
wire \branch_count_output[23]~42_combout ;
wire \pc_count_four_output[24]~45 ;
wire \pc_count_four_output[24]~44_combout ;
wire \pc_count_four_output[25]~47 ;
wire \pc_count_four_output[25]~46_combout ;
wire \branch_count_output[24]~45 ;
wire \branch_count_output[24]~44_combout ;
wire \branch_count_output[25]~47 ;
wire \branch_count_output[25]~46_combout ;
wire \branch_count_output[26]~49 ;
wire \branch_count_output[26]~48_combout ;
wire \pc_count_four_output[26]~49 ;
wire \pc_count_four_output[26]~48_combout ;
wire \pc_count_four_output[27]~51 ;
wire \pc_count_four_output[27]~50_combout ;
wire \pc_count_four_output[28]~53 ;
wire \pc_count_four_output[28]~52_combout ;
wire \branch_count_output[27]~51 ;
wire \branch_count_output[27]~50_combout ;
wire \pc_count_four_output[29]~55 ;
wire \pc_count_four_output[29]~54_combout ;
wire \branch_count_output[28]~53 ;
wire \branch_count_output[28]~52_combout ;
wire \branch_count_output[29]~55 ;
wire \branch_count_output[29]~54_combout ;
wire \pc_count_four_output[30]~57 ;
wire \pc_count_four_output[30]~56_combout ;
wire \pc_count_four_output[31]~58_combout ;
wire \branch_count_output[30]~57 ;
wire \branch_count_output[30]~56_combout ;
wire \branch_count_output[31]~58_combout ;
wire \IDEX|temp_halt_out_output~q ;
wire \EXMEM|temp_halt_out~q ;
wire \alusourceMUX|Mux30~0_combout ;
wire \EXMEM|temp_regwrite~q ;
wire \FORWADUNIT|always0~7_combout ;
wire \MEMWB|temp_regwrite~q ;
wire \FORWADUNIT|always0~8_combout ;
wire \FORWADUNIT|always0~12_combout ;
wire \ALUBMUX|alu_b_mux_output[1]~0_combout ;
wire \MEMTOREG|Mux30~1_combout ;
wire \FORWADUNIT|always0~13_combout ;
wire \FORWADUNIT|forwardb[1]~0_combout ;
wire \ALUBMUX|alu_b_mux_output[1]~1_combout ;
wire \alusourceMUX|Mux16~0_combout ;
wire \alusourceMUX|Mux30~1_combout ;
wire \FORWADUNIT|forwarda[1]~3_combout ;
wire \ALUAMUX|alu_a_mux_output[1]~1_combout ;
wire \MEMTOREG|Mux31~1_combout ;
wire \ALUBMUX|alu_b_mux_output[0]~2_combout ;
wire \alusourceMUX|Mux31~0_combout ;
wire \ALUBMUX|alu_b_mux_output[0]~3_combout ;
wire \ALUAMUX|alu_a_mux_output[0]~3_combout ;
wire \MEMTOREG|Mux29~1_combout ;
wire \ALUAMUX|alu_a_mux_output[2]~5_combout ;
wire \alusourceMUX|Mux31~1_combout ;
wire \MEMTOREG|Mux27~1_combout ;
wire \ALUAMUX|alu_a_mux_output[4]~7_combout ;
wire \MEMTOREG|Mux28~1_combout ;
wire \ALUAMUX|alu_a_mux_output[3]~8_combout ;
wire \ALUAMUX|alu_a_mux_output[3]~9_combout ;
wire \alusourceMUX|Mux29~0_combout ;
wire \ALUBMUX|alu_b_mux_output[2]~5_combout ;
wire \alusourceMUX|Mux29~1_combout ;
wire \MEMTOREG|Mux23~1_combout ;
wire \ALUAMUX|alu_a_mux_output[8]~11_combout ;
wire \MEMTOREG|Mux24~1_combout ;
wire \ALUAMUX|alu_a_mux_output[7]~13_combout ;
wire \MEMTOREG|Mux25~1_combout ;
wire \ALUAMUX|alu_a_mux_output[6]~15_combout ;
wire \MEMTOREG|Mux26~1_combout ;
wire \ALUAMUX|alu_a_mux_output[5]~17_combout ;
wire \alusourceMUX|Mux28~0_combout ;
wire \ALUBMUX|alu_b_mux_output[3]~7_combout ;
wire \alusourceMUX|Mux28~1_combout ;
wire \FORWADUNIT|always0~16_combout ;
wire \FORWADUNIT|always0~17_combout ;
wire \MEMTOREG|Mux15~1_combout ;
wire \ALUAMUX|alu_a_mux_output[16]~20_combout ;
wire \MEMTOREG|Mux17~1_combout ;
wire \ALUAMUX|alu_a_mux_output[14]~22_combout ;
wire \MEMTOREG|Mux16~1_combout ;
wire \ALUAMUX|alu_a_mux_output[15]~24_combout ;
wire \MEMTOREG|Mux18~1_combout ;
wire \ALUAMUX|alu_a_mux_output[13]~26_combout ;
wire \MEMTOREG|Mux19~1_combout ;
wire \ALUAMUX|alu_a_mux_output[12]~28_combout ;
wire \MEMTOREG|Mux21~1_combout ;
wire \ALUAMUX|alu_a_mux_output[10]~30_combout ;
wire \MEMTOREG|Mux20~1_combout ;
wire \ALUAMUX|alu_a_mux_output[11]~32_combout ;
wire \MEMTOREG|Mux22~1_combout ;
wire \ALUAMUX|alu_a_mux_output[9]~34_combout ;
wire \alusourceMUX|Mux27~0_combout ;
wire \ALUBMUX|alu_b_mux_output[4]~9_combout ;
wire \alusourceMUX|Mux27~1_combout ;
wire \MEMTOREG|Mux0~1_combout ;
wire \ALUAMUX|alu_a_mux_output[31]~36_combout ;
wire \MEMTOREG|Mux1~1_combout ;
wire \ALUAMUX|alu_a_mux_output[30]~38_combout ;
wire \MEMTOREG|Mux2~1_combout ;
wire \ALUAMUX|alu_a_mux_output[29]~40_combout ;
wire \MEMTOREG|Mux5~1_combout ;
wire \ALUAMUX|alu_a_mux_output[26]~42_combout ;
wire \MEMTOREG|Mux6~1_combout ;
wire \ALUAMUX|alu_a_mux_output[25]~44_combout ;
wire \MEMTOREG|Mux3~1_combout ;
wire \ALUAMUX|alu_a_mux_output[28]~46_combout ;
wire \MEMTOREG|Mux4~1_combout ;
wire \ALUAMUX|alu_a_mux_output[27]~48_combout ;
wire \MEMTOREG|Mux14~1_combout ;
wire \ALUAMUX|alu_a_mux_output[17]~50_combout ;
wire \MEMTOREG|Mux11~1_combout ;
wire \ALUAMUX|alu_a_mux_output[20]~52_combout ;
wire \MEMTOREG|Mux12~1_combout ;
wire \ALUAMUX|alu_a_mux_output[19]~54_combout ;
wire \MEMTOREG|Mux13~1_combout ;
wire \ALUAMUX|alu_a_mux_output[18]~56_combout ;
wire \MEMTOREG|Mux7~1_combout ;
wire \ALUAMUX|alu_a_mux_output[24]~58_combout ;
wire \MEMTOREG|Mux8~1_combout ;
wire \ALUAMUX|alu_a_mux_output[23]~60_combout ;
wire \MEMTOREG|Mux9~1_combout ;
wire \ALUAMUX|alu_a_mux_output[22]~62_combout ;
wire \MEMTOREG|Mux10~1_combout ;
wire \ALUAMUX|alu_a_mux_output[21]~64_combout ;
wire \ALUBMUX|alu_b_mux_output[15]~11_combout ;
wire \alusourceMUX|Mux16~1_combout ;
wire \ALUBMUX|alu_b_mux_output[12]~13_combout ;
wire \alusourceMUX|Mux19~0_combout ;
wire \ALUBMUX|alu_b_mux_output[27]~16_combout ;
wire \alusourceMUX|Mux4~0_combout ;
wire \ALUBMUX|alu_b_mux_output[18]~18_combout ;
wire \alusourceMUX|Mux13~0_combout ;
wire \ALUBMUX|alu_b_mux_output[17]~20_combout ;
wire \alusourceMUX|Mux14~0_combout ;
wire \ALUBMUX|alu_b_mux_output[16]~22_combout ;
wire \alusourceMUX|Mux15~0_combout ;
wire \ALUBMUX|alu_b_mux_output[31]~24_combout ;
wire \alusourceMUX|Mux0~0_combout ;
wire \ALUBMUX|alu_b_mux_output[30]~26_combout ;
wire \alusourceMUX|Mux1~0_combout ;
wire \ALUBMUX|alu_b_mux_output[29]~28_combout ;
wire \alusourceMUX|Mux2~0_combout ;
wire \ALUBMUX|alu_b_mux_output[28]~30_combout ;
wire \alusourceMUX|Mux3~0_combout ;
wire \ALUBMUX|alu_b_mux_output[26]~32_combout ;
wire \alusourceMUX|Mux5~0_combout ;
wire \ALUBMUX|alu_b_mux_output[25]~34_combout ;
wire \alusourceMUX|Mux6~0_combout ;
wire \ALUBMUX|alu_b_mux_output[24]~36_combout ;
wire \alusourceMUX|Mux7~0_combout ;
wire \ALUBMUX|alu_b_mux_output[23]~38_combout ;
wire \alusourceMUX|Mux8~0_combout ;
wire \ALUBMUX|alu_b_mux_output[22]~40_combout ;
wire \alusourceMUX|Mux9~0_combout ;
wire \ALUBMUX|alu_b_mux_output[21]~42_combout ;
wire \alusourceMUX|Mux10~0_combout ;
wire \ALUBMUX|alu_b_mux_output[20]~44_combout ;
wire \alusourceMUX|Mux11~0_combout ;
wire \ALUBMUX|alu_b_mux_output[19]~46_combout ;
wire \alusourceMUX|Mux12~0_combout ;
wire \alusourceMUX|Mux17~0_combout ;
wire \ALUBMUX|alu_b_mux_output[10]~48_combout ;
wire \alusourceMUX|Mux21~0_combout ;
wire \ALUBMUX|alu_b_mux_output[14]~50_combout ;
wire \ALUBMUX|alu_b_mux_output[9]~52_combout ;
wire \alusourceMUX|Mux22~0_combout ;
wire \ALUBMUX|alu_b_mux_output[8]~54_combout ;
wire \alusourceMUX|Mux23~0_combout ;
wire \ALUBMUX|alu_b_mux_output[7]~56_combout ;
wire \alusourceMUX|Mux24~0_combout ;
wire \ALUBMUX|alu_b_mux_output[6]~58_combout ;
wire \alusourceMUX|Mux25~0_combout ;
wire \ALUBMUX|alu_b_mux_output[5]~60_combout ;
wire \alusourceMUX|Mux26~0_combout ;
wire \ALUBMUX|alu_b_mux_output[13]~62_combout ;
wire \alusourceMUX|Mux18~0_combout ;
wire \ALUBMUX|alu_b_mux_output[11]~64_combout ;
wire \alusourceMUX|Mux20~0_combout ;
wire \ALU|Mux30~4_combout ;
wire \HAZARDUNIT|ex_mem_flush~0_combout ;
wire \HAZARDUNIT|ex_mem_flush~3_combout ;
wire \EXMEM|temp_branchSelect~q ;
wire \HAZARDUNIT|ex_mem_flush~4_combout ;
wire \HAZARDUNIT|ex_mem_flush~5_combout ;
wire \HAZARDUNIT|id_ex_wen~0_combout ;
wire \NPCMUX|Mux30~1_combout ;
wire \IDEX|temp_request_dmemREN_output~q ;
wire \HAZARDUNIT|use_after_load~6_combout ;
wire \HAZARDUNIT|pc_wen~2_combout ;
wire \IDEX|temp_request_dmemWEN_output~q ;
wire \alusourceMUX|Mux17~1_combout ;
wire \ALU|Mux31~9_combout ;
wire \NPCMUX|Mux31~2_combout ;
wire \ALU|Mux29~12_combout ;
wire \NPCMUX|Mux29~1_combout ;
wire \ALU|Mux28~6_combout ;
wire \NPCMUX|Mux28~1_combout ;
wire \ALUAMUX|alu_a_mux_output[3]~65_combout ;
wire \ALU|Mux26~6_combout ;
wire \NPCMUX|Mux26~1_combout ;
wire \ALU|Mux27~11_combout ;
wire \NPCMUX|Mux27~1_combout ;
wire \ALU|Mux24~6_combout ;
wire \NPCMUX|Mux24~1_combout ;
wire \ALU|Mux25~6_combout ;
wire \NPCMUX|Mux25~1_combout ;
wire \ALU|Mux22~0_combout ;
wire \ALU|Mux22~5_combout ;
wire \ALU|Mux19~6_combout ;
wire \NPCMUX|Mux22~1_combout ;
wire \ALU|Mux23~0_combout ;
wire \ALU|Mux23~5_combout ;
wire \NPCMUX|Mux23~1_combout ;
wire \ALU|Mux20~0_combout ;
wire \ALU|Mux20~5_combout ;
wire \NPCMUX|Mux20~1_combout ;
wire \ALU|Mux21~0_combout ;
wire \ALU|Mux21~5_combout ;
wire \NPCMUX|Mux21~1_combout ;
wire \ALU|Mux18~0_combout ;
wire \ALU|Mux18~5_combout ;
wire \NPCMUX|Mux18~1_combout ;
wire \ALU|Mux19~7_combout ;
wire \ALU|Mux19~12_combout ;
wire \NPCMUX|Mux19~1_combout ;
wire \ALU|Mux16~0_combout ;
wire \ALU|Mux16~5_combout ;
wire \NPCMUX|Mux16~1_combout ;
wire \ALU|Mux17~0_combout ;
wire \ALU|Mux17~5_combout ;
wire \NPCMUX|Mux17~1_combout ;
wire \ALU|Mux14~0_combout ;
wire \ALU|Mux14~4_combout ;
wire \NPCMUX|Mux14~1_combout ;
wire \ALU|Mux15~0_combout ;
wire \ALU|Mux15~4_combout ;
wire \NPCMUX|Mux15~1_combout ;
wire \ALU|Mux12~3_combout ;
wire \ALU|Mux12~8_combout ;
wire \NPCMUX|Mux12~1_combout ;
wire \ALU|Mux13~0_combout ;
wire \ALU|Mux13~5_combout ;
wire \NPCMUX|Mux13~1_combout ;
wire \ALU|Mux11~0_combout ;
wire \ALU|Mux11~5_combout ;
wire \NPCMUX|Mux11~1_combout ;
wire \ALU|Mux10~0_combout ;
wire \ALU|Mux10~5_combout ;
wire \NPCMUX|Mux10~1_combout ;
wire \ALU|Mux8~0_combout ;
wire \ALU|Mux8~5_combout ;
wire \NPCMUX|Mux8~1_combout ;
wire \ALU|Mux9~0_combout ;
wire \ALU|Mux9~5_combout ;
wire \NPCMUX|Mux9~1_combout ;
wire \ALU|Mux6~7_combout ;
wire \NPCMUX|Mux6~1_combout ;
wire \NPCMUX|Mux7~1_combout ;
wire \NPCMUX|Mux5~1_combout ;
wire \ALU|Mux4~7_combout ;
wire \NPCMUX|Mux4~1_combout ;
wire \ALU|Mux2~14_combout ;
wire \NPCMUX|Mux2~1_combout ;
wire \ALU|Mux3~9_combout ;
wire \NPCMUX|Mux3~3_combout ;
wire \ALU|Mux0~0_combout ;
wire \ALU|Mux0~7_combout ;
wire \NPCMUX|Mux0~1_combout ;
wire \ALU|Mux1~2_combout ;
wire \NPCMUX|Mux1~1_combout ;
wire \CONTROLUNIT|Equal3~0_combout ;
wire \IDEX|temp_branch_output~0_combout ;
wire \CONTROLUNIT|Equal3~1_combout ;
wire \CONTROLUNIT|Equal3~9_combout ;
wire \EXTENDER|extended_imm[16]~0_combout ;
wire \CONTROLUNIT|WideOr8~0_combout ;
wire \CONTROLUNIT|WideOr2~0_combout ;
wire \HAZARDUNIT|id_ex_flush~combout ;
wire \CONTROLUNIT|WideOr4~0_combout ;
wire \IDEX|temp_ALUsrc_output~3_combout ;
wire \REGISTER|Mux62~9_combout ;
wire \REGISTER|Mux62~19_combout ;
wire \IDEX|temp_regwrite_output~q ;
wire \REGISTER|Mux30~9_combout ;
wire \REGISTER|Mux30~19_combout ;
wire \CONTROLUNIT|WideOr7~0_combout ;
wire \CONTROLUNIT|WideOr1~0_combout ;
wire \REGISTER|Mux63~9_combout ;
wire \REGISTER|Mux63~19_combout ;
wire \REGISTER|Mux31~9_combout ;
wire \REGISTER|Mux31~19_combout ;
wire \REGISTER|Mux29~9_combout ;
wire \REGISTER|Mux29~19_combout ;
wire \REGISTER|Mux27~9_combout ;
wire \REGISTER|Mux27~19_combout ;
wire \REGISTER|Mux28~9_combout ;
wire \REGISTER|Mux28~19_combout ;
wire \REGISTER|Mux61~9_combout ;
wire \REGISTER|Mux61~19_combout ;
wire \REGISTER|Mux23~9_combout ;
wire \REGISTER|Mux23~19_combout ;
wire \REGISTER|Mux24~9_combout ;
wire \REGISTER|Mux24~19_combout ;
wire \REGISTER|Mux25~9_combout ;
wire \REGISTER|Mux25~19_combout ;
wire \REGISTER|Mux26~9_combout ;
wire \REGISTER|Mux26~19_combout ;
wire \REGISTER|Mux60~9_combout ;
wire \REGISTER|Mux60~19_combout ;
wire \REGISTER|Mux15~9_combout ;
wire \REGISTER|Mux15~19_combout ;
wire \REGISTER|Mux17~9_combout ;
wire \REGISTER|Mux17~19_combout ;
wire \REGISTER|Mux16~9_combout ;
wire \REGISTER|Mux16~19_combout ;
wire \REGISTER|Mux18~9_combout ;
wire \REGISTER|Mux18~19_combout ;
wire \REGISTER|Mux19~9_combout ;
wire \REGISTER|Mux19~19_combout ;
wire \REGISTER|Mux21~9_combout ;
wire \REGISTER|Mux21~19_combout ;
wire \REGISTER|Mux20~9_combout ;
wire \REGISTER|Mux20~19_combout ;
wire \REGISTER|Mux22~9_combout ;
wire \REGISTER|Mux22~19_combout ;
wire \REGISTER|Mux59~9_combout ;
wire \REGISTER|Mux59~19_combout ;
wire \REGISTER|Mux0~9_combout ;
wire \REGISTER|Mux0~19_combout ;
wire \REGISTER|Mux1~9_combout ;
wire \REGISTER|Mux1~19_combout ;
wire \REGISTER|Mux2~9_combout ;
wire \REGISTER|Mux2~19_combout ;
wire \REGISTER|Mux5~9_combout ;
wire \REGISTER|Mux5~19_combout ;
wire \REGISTER|Mux6~9_combout ;
wire \REGISTER|Mux6~19_combout ;
wire \REGISTER|Mux3~9_combout ;
wire \REGISTER|Mux3~19_combout ;
wire \REGISTER|Mux4~9_combout ;
wire \REGISTER|Mux4~19_combout ;
wire \REGISTER|Mux14~9_combout ;
wire \REGISTER|Mux14~19_combout ;
wire \REGISTER|Mux11~9_combout ;
wire \REGISTER|Mux11~19_combout ;
wire \REGISTER|Mux12~9_combout ;
wire \REGISTER|Mux12~19_combout ;
wire \REGISTER|Mux13~9_combout ;
wire \REGISTER|Mux13~19_combout ;
wire \REGISTER|Mux7~9_combout ;
wire \REGISTER|Mux7~19_combout ;
wire \REGISTER|Mux8~9_combout ;
wire \REGISTER|Mux8~19_combout ;
wire \REGISTER|Mux9~9_combout ;
wire \REGISTER|Mux9~19_combout ;
wire \REGISTER|Mux10~9_combout ;
wire \REGISTER|Mux10~19_combout ;
wire \REGISTER|Mux48~9_combout ;
wire \REGISTER|Mux48~19_combout ;
wire \REGISTER|Mux51~9_combout ;
wire \REGISTER|Mux51~19_combout ;
wire \REGISTER|Mux36~9_combout ;
wire \REGISTER|Mux36~19_combout ;
wire \CONTROLUNIT|WideOr5~0_combout ;
wire \EXTENDER|extended_imm[16]~2_combout ;
wire \REGISTER|Mux45~9_combout ;
wire \REGISTER|Mux45~19_combout ;
wire \REGISTER|Mux46~9_combout ;
wire \REGISTER|Mux46~19_combout ;
wire \REGISTER|Mux47~9_combout ;
wire \REGISTER|Mux47~19_combout ;
wire \REGISTER|Mux32~9_combout ;
wire \REGISTER|Mux32~19_combout ;
wire \REGISTER|Mux33~9_combout ;
wire \REGISTER|Mux33~19_combout ;
wire \REGISTER|Mux34~9_combout ;
wire \REGISTER|Mux34~19_combout ;
wire \REGISTER|Mux35~9_combout ;
wire \REGISTER|Mux35~19_combout ;
wire \REGISTER|Mux37~9_combout ;
wire \REGISTER|Mux37~19_combout ;
wire \REGISTER|Mux38~9_combout ;
wire \REGISTER|Mux38~19_combout ;
wire \REGISTER|Mux39~9_combout ;
wire \REGISTER|Mux39~19_combout ;
wire \REGISTER|Mux40~9_combout ;
wire \REGISTER|Mux40~19_combout ;
wire \REGISTER|Mux41~9_combout ;
wire \REGISTER|Mux41~19_combout ;
wire \REGISTER|Mux42~9_combout ;
wire \REGISTER|Mux42~19_combout ;
wire \REGISTER|Mux43~9_combout ;
wire \REGISTER|Mux43~19_combout ;
wire \REGISTER|Mux44~9_combout ;
wire \REGISTER|Mux44~19_combout ;
wire \REGISTER|Mux53~9_combout ;
wire \REGISTER|Mux53~19_combout ;
wire \REGISTER|Mux49~9_combout ;
wire \REGISTER|Mux49~19_combout ;
wire \REGISTER|Mux54~9_combout ;
wire \REGISTER|Mux54~19_combout ;
wire \REGISTER|Mux55~9_combout ;
wire \REGISTER|Mux55~19_combout ;
wire \REGISTER|Mux56~9_combout ;
wire \REGISTER|Mux56~19_combout ;
wire \REGISTER|Mux57~9_combout ;
wire \REGISTER|Mux57~19_combout ;
wire \REGISTER|Mux58~9_combout ;
wire \REGISTER|Mux58~19_combout ;
wire \REGISTER|Mux50~9_combout ;
wire \REGISTER|Mux50~19_combout ;
wire \REGISTER|Mux52~9_combout ;
wire \REGISTER|Mux52~19_combout ;
wire \CONTROLUNIT|WideOr6~0_combout ;
wire \CONTROLUNIT|WideOr0~0_combout ;
wire \CONTROLUNIT|halt_out~0_combout ;
wire \IDEX|temp_branch_output~q ;
wire \ALU|Equal0~22_combout ;
wire \HAZARDUNIT|pc_wen~3_combout ;
wire \CONTROLUNIT|halt_out~3_combout ;
wire \CONTROLUNIT|WideOr3~0_combout ;
wire \CONTROLUNIT|WideOr10~0_combout ;
wire \CONTROLUNIT|memtoreg~0_combout ;
wire \CONTROLUNIT|WideOr9~0_combout ;
wire \FORWADUNIT|always0~18_combout ;
wire \FORWADUNIT|always0~19_combout ;
wire \ALU|Mux1~10_combout ;
wire \ALU|Mux5~8_combout ;
wire \ALU|Mux7~7_combout ;
wire [31:0] \IFID|temp_imemload_output ;
wire [31:0] \IFID|temp_NPC_output ;
wire [31:0] \IDEX|temp_signzerovalue_output ;
wire [1:0] \IDEX|temp_regdst_output ;
wire [31:0] \IDEX|temp_rdat_two_output ;
wire [31:0] \IDEX|temp_rdat_one_output ;
wire [2:0] \IDEX|temp_pcselect_output ;
wire [1:0] \IDEX|temp_memtoreg_output ;
wire [31:0] \IDEX|temp_imemload_output ;
wire [31:0] \IDEX|temp_NPC_output ;
wire [1:0] \IDEX|temp_ALUsrc_output ;
wire [3:0] \IDEX|temp_ALUop_output ;
wire [31:0] \EXMEM|temp_signZero ;
wire [31:0] \EXMEM|temp_rdat1 ;
wire [1:0] \EXMEM|temp_pcselect ;
wire [31:0] \EXMEM|temp_npc ;
wire [1:0] \EXMEM|temp_memtoreg ;
wire [31:0] \EXMEM|temp_iMemLoad ;
wire [4:0] \EXMEM|temp_branchDest ;
wire [31:0] \MEMWB|temp_upper16 ;
wire [31:0] \MEMWB|temp_npc ;
wire [1:0] \MEMWB|temp_memtoreg ;
wire [31:0] \MEMWB|temp_dMemLoad ;
wire [4:0] \MEMWB|temp_branchDest ;
wire [31:0] \MEMWB|temp_aluResult ;


alu_b_mux ALUBMUX(
	.temp_aluResult_1(temp_aluResult_1),
	.temp_aluResult_0(temp_aluResult_0),
	.temp_aluResult_2(temp_aluResult_2),
	.temp_aluResult_3(temp_aluResult_3),
	.temp_aluResult_5(temp_aluResult_5),
	.temp_aluResult_4(temp_aluResult_4),
	.temp_aluResult_7(temp_aluResult_7),
	.temp_aluResult_6(temp_aluResult_6),
	.temp_aluResult_9(temp_aluResult_9),
	.temp_aluResult_8(temp_aluResult_8),
	.temp_aluResult_11(temp_aluResult_11),
	.temp_aluResult_10(temp_aluResult_10),
	.temp_aluResult_13(temp_aluResult_13),
	.temp_aluResult_12(temp_aluResult_12),
	.temp_aluResult_15(temp_aluResult_15),
	.temp_aluResult_14(temp_aluResult_14),
	.temp_aluResult_17(temp_aluResult_17),
	.temp_aluResult_16(temp_aluResult_16),
	.temp_aluResult_19(temp_aluResult_19),
	.temp_aluResult_18(temp_aluResult_18),
	.temp_aluResult_20(temp_aluResult_20),
	.temp_aluResult_21(temp_aluResult_21),
	.temp_aluResult_23(temp_aluResult_23),
	.temp_aluResult_22(temp_aluResult_22),
	.temp_aluResult_25(temp_aluResult_25),
	.temp_aluResult_24(temp_aluResult_24),
	.temp_aluResult_26(temp_aluResult_26),
	.temp_aluResult_27(temp_aluResult_27),
	.temp_aluResult_29(temp_aluResult_29),
	.temp_aluResult_28(temp_aluResult_28),
	.temp_aluResult_31(temp_aluResult_31),
	.temp_aluResult_30(temp_aluResult_30),
	.temp_rdat_two_output_1(\IDEX|temp_rdat_two_output [1]),
	.always0(\FORWADUNIT|always0~7_combout ),
	.always01(\FORWADUNIT|always0~8_combout ),
	.always02(\FORWADUNIT|always0~12_combout ),
	.alu_b_mux_output_1(\ALUBMUX|alu_b_mux_output[1]~0_combout ),
	.Mux30(\MEMTOREG|Mux30~1_combout ),
	.always03(\FORWADUNIT|always0~13_combout ),
	.forwardb_1(\FORWADUNIT|forwardb[1]~0_combout ),
	.alu_b_mux_output_11(\ALUBMUX|alu_b_mux_output[1]~1_combout ),
	.Mux31(\MEMTOREG|Mux31~1_combout ),
	.alu_b_mux_output_0(\ALUBMUX|alu_b_mux_output[0]~2_combout ),
	.temp_rdat_two_output_0(\IDEX|temp_rdat_two_output [0]),
	.alu_b_mux_output_01(\ALUBMUX|alu_b_mux_output[0]~3_combout ),
	.Mux29(\MEMTOREG|Mux29~1_combout ),
	.Mux27(\MEMTOREG|Mux27~1_combout ),
	.Mux28(\MEMTOREG|Mux28~1_combout ),
	.temp_rdat_two_output_2(\IDEX|temp_rdat_two_output [2]),
	.alu_b_mux_output_2(\ALUBMUX|alu_b_mux_output[2]~5_combout ),
	.Mux23(\MEMTOREG|Mux23~1_combout ),
	.Mux24(\MEMTOREG|Mux24~1_combout ),
	.Mux25(\MEMTOREG|Mux25~1_combout ),
	.Mux26(\MEMTOREG|Mux26~1_combout ),
	.temp_rdat_two_output_3(\IDEX|temp_rdat_two_output [3]),
	.alu_b_mux_output_3(\ALUBMUX|alu_b_mux_output[3]~7_combout ),
	.Mux15(\MEMTOREG|Mux15~1_combout ),
	.temp_iMemLoad_0(\EXMEM|temp_iMemLoad [0]),
	.Mux17(\MEMTOREG|Mux17~1_combout ),
	.Mux16(\MEMTOREG|Mux16~1_combout ),
	.Mux18(\MEMTOREG|Mux18~1_combout ),
	.Mux19(\MEMTOREG|Mux19~1_combout ),
	.Mux21(\MEMTOREG|Mux21~1_combout ),
	.Mux20(\MEMTOREG|Mux20~1_combout ),
	.Mux22(\MEMTOREG|Mux22~1_combout ),
	.temp_rdat_two_output_4(\IDEX|temp_rdat_two_output [4]),
	.alu_b_mux_output_4(\ALUBMUX|alu_b_mux_output[4]~9_combout ),
	.Mux0(\MEMTOREG|Mux0~1_combout ),
	.temp_iMemLoad_15(\EXMEM|temp_iMemLoad [15]),
	.Mux1(\MEMTOREG|Mux1~1_combout ),
	.temp_iMemLoad_14(\EXMEM|temp_iMemLoad [14]),
	.Mux2(\MEMTOREG|Mux2~1_combout ),
	.temp_iMemLoad_13(\EXMEM|temp_iMemLoad [13]),
	.Mux5(\MEMTOREG|Mux5~1_combout ),
	.temp_iMemLoad_10(\EXMEM|temp_iMemLoad [10]),
	.Mux6(\MEMTOREG|Mux6~1_combout ),
	.temp_iMemLoad_9(\EXMEM|temp_iMemLoad [9]),
	.Mux3(\MEMTOREG|Mux3~1_combout ),
	.temp_iMemLoad_12(\EXMEM|temp_iMemLoad [12]),
	.Mux4(\MEMTOREG|Mux4~1_combout ),
	.temp_iMemLoad_11(\EXMEM|temp_iMemLoad [11]),
	.Mux14(\MEMTOREG|Mux14~1_combout ),
	.temp_iMemLoad_1(\EXMEM|temp_iMemLoad [1]),
	.Mux11(\MEMTOREG|Mux11~1_combout ),
	.temp_iMemLoad_4(\EXMEM|temp_iMemLoad [4]),
	.Mux12(\MEMTOREG|Mux12~1_combout ),
	.temp_iMemLoad_3(\EXMEM|temp_iMemLoad [3]),
	.Mux13(\MEMTOREG|Mux13~1_combout ),
	.temp_iMemLoad_2(\EXMEM|temp_iMemLoad [2]),
	.Mux7(\MEMTOREG|Mux7~1_combout ),
	.temp_iMemLoad_8(\EXMEM|temp_iMemLoad [8]),
	.Mux8(\MEMTOREG|Mux8~1_combout ),
	.temp_iMemLoad_7(\EXMEM|temp_iMemLoad [7]),
	.Mux9(\MEMTOREG|Mux9~1_combout ),
	.temp_iMemLoad_6(\EXMEM|temp_iMemLoad [6]),
	.Mux10(\MEMTOREG|Mux10~1_combout ),
	.temp_iMemLoad_5(\EXMEM|temp_iMemLoad [5]),
	.temp_rdat_two_output_15(\IDEX|temp_rdat_two_output [15]),
	.alu_b_mux_output_15(\ALUBMUX|alu_b_mux_output[15]~11_combout ),
	.temp_rdat_two_output_12(\IDEX|temp_rdat_two_output [12]),
	.alu_b_mux_output_12(\ALUBMUX|alu_b_mux_output[12]~13_combout ),
	.temp_rdat_two_output_27(\IDEX|temp_rdat_two_output [27]),
	.alu_b_mux_output_27(\ALUBMUX|alu_b_mux_output[27]~16_combout ),
	.temp_rdat_two_output_18(\IDEX|temp_rdat_two_output [18]),
	.alu_b_mux_output_18(\ALUBMUX|alu_b_mux_output[18]~18_combout ),
	.temp_rdat_two_output_17(\IDEX|temp_rdat_two_output [17]),
	.alu_b_mux_output_17(\ALUBMUX|alu_b_mux_output[17]~20_combout ),
	.temp_rdat_two_output_16(\IDEX|temp_rdat_two_output [16]),
	.alu_b_mux_output_16(\ALUBMUX|alu_b_mux_output[16]~22_combout ),
	.temp_rdat_two_output_31(\IDEX|temp_rdat_two_output [31]),
	.alu_b_mux_output_31(\ALUBMUX|alu_b_mux_output[31]~24_combout ),
	.temp_rdat_two_output_30(\IDEX|temp_rdat_two_output [30]),
	.alu_b_mux_output_30(\ALUBMUX|alu_b_mux_output[30]~26_combout ),
	.temp_rdat_two_output_29(\IDEX|temp_rdat_two_output [29]),
	.alu_b_mux_output_29(\ALUBMUX|alu_b_mux_output[29]~28_combout ),
	.temp_rdat_two_output_28(\IDEX|temp_rdat_two_output [28]),
	.alu_b_mux_output_28(\ALUBMUX|alu_b_mux_output[28]~30_combout ),
	.temp_rdat_two_output_26(\IDEX|temp_rdat_two_output [26]),
	.alu_b_mux_output_26(\ALUBMUX|alu_b_mux_output[26]~32_combout ),
	.temp_rdat_two_output_25(\IDEX|temp_rdat_two_output [25]),
	.alu_b_mux_output_25(\ALUBMUX|alu_b_mux_output[25]~34_combout ),
	.temp_rdat_two_output_24(\IDEX|temp_rdat_two_output [24]),
	.alu_b_mux_output_24(\ALUBMUX|alu_b_mux_output[24]~36_combout ),
	.temp_rdat_two_output_23(\IDEX|temp_rdat_two_output [23]),
	.alu_b_mux_output_23(\ALUBMUX|alu_b_mux_output[23]~38_combout ),
	.temp_rdat_two_output_22(\IDEX|temp_rdat_two_output [22]),
	.alu_b_mux_output_22(\ALUBMUX|alu_b_mux_output[22]~40_combout ),
	.temp_rdat_two_output_21(\IDEX|temp_rdat_two_output [21]),
	.alu_b_mux_output_21(\ALUBMUX|alu_b_mux_output[21]~42_combout ),
	.temp_rdat_two_output_20(\IDEX|temp_rdat_two_output [20]),
	.alu_b_mux_output_20(\ALUBMUX|alu_b_mux_output[20]~44_combout ),
	.temp_rdat_two_output_19(\IDEX|temp_rdat_two_output [19]),
	.alu_b_mux_output_19(\ALUBMUX|alu_b_mux_output[19]~46_combout ),
	.temp_rdat_two_output_10(\IDEX|temp_rdat_two_output [10]),
	.alu_b_mux_output_10(\ALUBMUX|alu_b_mux_output[10]~48_combout ),
	.temp_rdat_two_output_14(\IDEX|temp_rdat_two_output [14]),
	.alu_b_mux_output_14(\ALUBMUX|alu_b_mux_output[14]~50_combout ),
	.temp_rdat_two_output_9(\IDEX|temp_rdat_two_output [9]),
	.alu_b_mux_output_9(\ALUBMUX|alu_b_mux_output[9]~52_combout ),
	.temp_rdat_two_output_8(\IDEX|temp_rdat_two_output [8]),
	.alu_b_mux_output_8(\ALUBMUX|alu_b_mux_output[8]~54_combout ),
	.temp_rdat_two_output_7(\IDEX|temp_rdat_two_output [7]),
	.alu_b_mux_output_7(\ALUBMUX|alu_b_mux_output[7]~56_combout ),
	.temp_rdat_two_output_6(\IDEX|temp_rdat_two_output [6]),
	.alu_b_mux_output_6(\ALUBMUX|alu_b_mux_output[6]~58_combout ),
	.temp_rdat_two_output_5(\IDEX|temp_rdat_two_output [5]),
	.alu_b_mux_output_5(\ALUBMUX|alu_b_mux_output[5]~60_combout ),
	.temp_rdat_two_output_13(\IDEX|temp_rdat_two_output [13]),
	.alu_b_mux_output_13(\ALUBMUX|alu_b_mux_output[13]~62_combout ),
	.temp_rdat_two_output_11(\IDEX|temp_rdat_two_output [11]),
	.alu_b_mux_output_111(\ALUBMUX|alu_b_mux_output[11]~64_combout ),
	.always04(\FORWADUNIT|always0~18_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

alu_a_mux ALUAMUX(
	.temp_aluResult_1(temp_aluResult_1),
	.temp_aluResult_0(temp_aluResult_0),
	.temp_aluResult_2(temp_aluResult_2),
	.temp_aluResult_3(temp_aluResult_3),
	.temp_aluResult_5(temp_aluResult_5),
	.temp_aluResult_4(temp_aluResult_4),
	.temp_aluResult_7(temp_aluResult_7),
	.temp_aluResult_6(temp_aluResult_6),
	.temp_aluResult_9(temp_aluResult_9),
	.temp_aluResult_8(temp_aluResult_8),
	.temp_aluResult_11(temp_aluResult_11),
	.temp_aluResult_10(temp_aluResult_10),
	.temp_aluResult_13(temp_aluResult_13),
	.temp_aluResult_12(temp_aluResult_12),
	.temp_aluResult_15(temp_aluResult_15),
	.temp_aluResult_14(temp_aluResult_14),
	.temp_aluResult_17(temp_aluResult_17),
	.temp_aluResult_16(temp_aluResult_16),
	.temp_aluResult_19(temp_aluResult_19),
	.temp_aluResult_18(temp_aluResult_18),
	.temp_aluResult_20(temp_aluResult_20),
	.temp_aluResult_21(temp_aluResult_21),
	.temp_aluResult_23(temp_aluResult_23),
	.temp_aluResult_22(temp_aluResult_22),
	.temp_aluResult_25(temp_aluResult_25),
	.temp_aluResult_24(temp_aluResult_24),
	.temp_aluResult_26(temp_aluResult_26),
	.temp_aluResult_27(temp_aluResult_27),
	.temp_aluResult_29(temp_aluResult_29),
	.temp_aluResult_28(temp_aluResult_28),
	.temp_aluResult_31(temp_aluResult_31),
	.temp_aluResult_30(temp_aluResult_30),
	.always0(\FORWADUNIT|always0~8_combout ),
	.Mux30(\MEMTOREG|Mux30~1_combout ),
	.forwarda_1(\FORWADUNIT|forwarda[1]~3_combout ),
	.temp_rdat_one_output_1(\IDEX|temp_rdat_one_output [1]),
	.alu_a_mux_output_1(\ALUAMUX|alu_a_mux_output[1]~1_combout ),
	.Mux31(\MEMTOREG|Mux31~1_combout ),
	.temp_rdat_one_output_0(\IDEX|temp_rdat_one_output [0]),
	.alu_a_mux_output_0(\ALUAMUX|alu_a_mux_output[0]~3_combout ),
	.Mux29(\MEMTOREG|Mux29~1_combout ),
	.temp_rdat_one_output_2(\IDEX|temp_rdat_one_output [2]),
	.alu_a_mux_output_2(\ALUAMUX|alu_a_mux_output[2]~5_combout ),
	.Mux27(\MEMTOREG|Mux27~1_combout ),
	.temp_rdat_one_output_4(\IDEX|temp_rdat_one_output [4]),
	.alu_a_mux_output_4(\ALUAMUX|alu_a_mux_output[4]~7_combout ),
	.Mux28(\MEMTOREG|Mux28~1_combout ),
	.alu_a_mux_output_3(\ALUAMUX|alu_a_mux_output[3]~8_combout ),
	.temp_rdat_one_output_3(\IDEX|temp_rdat_one_output [3]),
	.alu_a_mux_output_31(\ALUAMUX|alu_a_mux_output[3]~9_combout ),
	.Mux23(\MEMTOREG|Mux23~1_combout ),
	.temp_rdat_one_output_8(\IDEX|temp_rdat_one_output [8]),
	.alu_a_mux_output_8(\ALUAMUX|alu_a_mux_output[8]~11_combout ),
	.Mux24(\MEMTOREG|Mux24~1_combout ),
	.temp_rdat_one_output_7(\IDEX|temp_rdat_one_output [7]),
	.alu_a_mux_output_7(\ALUAMUX|alu_a_mux_output[7]~13_combout ),
	.Mux25(\MEMTOREG|Mux25~1_combout ),
	.temp_rdat_one_output_6(\IDEX|temp_rdat_one_output [6]),
	.alu_a_mux_output_6(\ALUAMUX|alu_a_mux_output[6]~15_combout ),
	.Mux26(\MEMTOREG|Mux26~1_combout ),
	.temp_rdat_one_output_5(\IDEX|temp_rdat_one_output [5]),
	.alu_a_mux_output_5(\ALUAMUX|alu_a_mux_output[5]~17_combout ),
	.temp_rdat_one_output_16(\IDEX|temp_rdat_one_output [16]),
	.always01(\FORWADUNIT|always0~16_combout ),
	.always02(\FORWADUNIT|always0~17_combout ),
	.Mux15(\MEMTOREG|Mux15~1_combout ),
	.temp_iMemLoad_0(\EXMEM|temp_iMemLoad [0]),
	.alu_a_mux_output_16(\ALUAMUX|alu_a_mux_output[16]~20_combout ),
	.Mux17(\MEMTOREG|Mux17~1_combout ),
	.temp_rdat_one_output_14(\IDEX|temp_rdat_one_output [14]),
	.alu_a_mux_output_14(\ALUAMUX|alu_a_mux_output[14]~22_combout ),
	.Mux16(\MEMTOREG|Mux16~1_combout ),
	.temp_rdat_one_output_15(\IDEX|temp_rdat_one_output [15]),
	.alu_a_mux_output_15(\ALUAMUX|alu_a_mux_output[15]~24_combout ),
	.Mux18(\MEMTOREG|Mux18~1_combout ),
	.temp_rdat_one_output_13(\IDEX|temp_rdat_one_output [13]),
	.alu_a_mux_output_13(\ALUAMUX|alu_a_mux_output[13]~26_combout ),
	.Mux19(\MEMTOREG|Mux19~1_combout ),
	.temp_rdat_one_output_12(\IDEX|temp_rdat_one_output [12]),
	.alu_a_mux_output_12(\ALUAMUX|alu_a_mux_output[12]~28_combout ),
	.Mux21(\MEMTOREG|Mux21~1_combout ),
	.temp_rdat_one_output_10(\IDEX|temp_rdat_one_output [10]),
	.alu_a_mux_output_10(\ALUAMUX|alu_a_mux_output[10]~30_combout ),
	.Mux20(\MEMTOREG|Mux20~1_combout ),
	.temp_rdat_one_output_11(\IDEX|temp_rdat_one_output [11]),
	.alu_a_mux_output_11(\ALUAMUX|alu_a_mux_output[11]~32_combout ),
	.Mux22(\MEMTOREG|Mux22~1_combout ),
	.temp_rdat_one_output_9(\IDEX|temp_rdat_one_output [9]),
	.alu_a_mux_output_9(\ALUAMUX|alu_a_mux_output[9]~34_combout ),
	.temp_rdat_one_output_31(\IDEX|temp_rdat_one_output [31]),
	.Mux0(\MEMTOREG|Mux0~1_combout ),
	.temp_iMemLoad_15(\EXMEM|temp_iMemLoad [15]),
	.alu_a_mux_output_311(\ALUAMUX|alu_a_mux_output[31]~36_combout ),
	.temp_rdat_one_output_30(\IDEX|temp_rdat_one_output [30]),
	.Mux1(\MEMTOREG|Mux1~1_combout ),
	.temp_iMemLoad_14(\EXMEM|temp_iMemLoad [14]),
	.alu_a_mux_output_30(\ALUAMUX|alu_a_mux_output[30]~38_combout ),
	.temp_rdat_one_output_29(\IDEX|temp_rdat_one_output [29]),
	.Mux2(\MEMTOREG|Mux2~1_combout ),
	.temp_iMemLoad_13(\EXMEM|temp_iMemLoad [13]),
	.alu_a_mux_output_29(\ALUAMUX|alu_a_mux_output[29]~40_combout ),
	.temp_rdat_one_output_26(\IDEX|temp_rdat_one_output [26]),
	.Mux5(\MEMTOREG|Mux5~1_combout ),
	.temp_iMemLoad_10(\EXMEM|temp_iMemLoad [10]),
	.alu_a_mux_output_26(\ALUAMUX|alu_a_mux_output[26]~42_combout ),
	.temp_rdat_one_output_25(\IDEX|temp_rdat_one_output [25]),
	.Mux6(\MEMTOREG|Mux6~1_combout ),
	.temp_iMemLoad_9(\EXMEM|temp_iMemLoad [9]),
	.alu_a_mux_output_25(\ALUAMUX|alu_a_mux_output[25]~44_combout ),
	.temp_rdat_one_output_28(\IDEX|temp_rdat_one_output [28]),
	.Mux3(\MEMTOREG|Mux3~1_combout ),
	.temp_iMemLoad_12(\EXMEM|temp_iMemLoad [12]),
	.alu_a_mux_output_28(\ALUAMUX|alu_a_mux_output[28]~46_combout ),
	.temp_rdat_one_output_27(\IDEX|temp_rdat_one_output [27]),
	.Mux4(\MEMTOREG|Mux4~1_combout ),
	.temp_iMemLoad_11(\EXMEM|temp_iMemLoad [11]),
	.alu_a_mux_output_27(\ALUAMUX|alu_a_mux_output[27]~48_combout ),
	.temp_rdat_one_output_17(\IDEX|temp_rdat_one_output [17]),
	.Mux14(\MEMTOREG|Mux14~1_combout ),
	.temp_iMemLoad_1(\EXMEM|temp_iMemLoad [1]),
	.alu_a_mux_output_17(\ALUAMUX|alu_a_mux_output[17]~50_combout ),
	.temp_rdat_one_output_20(\IDEX|temp_rdat_one_output [20]),
	.Mux11(\MEMTOREG|Mux11~1_combout ),
	.temp_iMemLoad_4(\EXMEM|temp_iMemLoad [4]),
	.alu_a_mux_output_20(\ALUAMUX|alu_a_mux_output[20]~52_combout ),
	.temp_rdat_one_output_19(\IDEX|temp_rdat_one_output [19]),
	.Mux12(\MEMTOREG|Mux12~1_combout ),
	.temp_iMemLoad_3(\EXMEM|temp_iMemLoad [3]),
	.alu_a_mux_output_19(\ALUAMUX|alu_a_mux_output[19]~54_combout ),
	.temp_rdat_one_output_18(\IDEX|temp_rdat_one_output [18]),
	.Mux13(\MEMTOREG|Mux13~1_combout ),
	.temp_iMemLoad_2(\EXMEM|temp_iMemLoad [2]),
	.alu_a_mux_output_18(\ALUAMUX|alu_a_mux_output[18]~56_combout ),
	.temp_rdat_one_output_24(\IDEX|temp_rdat_one_output [24]),
	.Mux7(\MEMTOREG|Mux7~1_combout ),
	.temp_iMemLoad_8(\EXMEM|temp_iMemLoad [8]),
	.alu_a_mux_output_24(\ALUAMUX|alu_a_mux_output[24]~58_combout ),
	.temp_rdat_one_output_23(\IDEX|temp_rdat_one_output [23]),
	.Mux8(\MEMTOREG|Mux8~1_combout ),
	.temp_iMemLoad_7(\EXMEM|temp_iMemLoad [7]),
	.alu_a_mux_output_23(\ALUAMUX|alu_a_mux_output[23]~60_combout ),
	.temp_rdat_one_output_22(\IDEX|temp_rdat_one_output [22]),
	.Mux9(\MEMTOREG|Mux9~1_combout ),
	.temp_iMemLoad_6(\EXMEM|temp_iMemLoad [6]),
	.alu_a_mux_output_22(\ALUAMUX|alu_a_mux_output[22]~62_combout ),
	.temp_rdat_one_output_21(\IDEX|temp_rdat_one_output [21]),
	.Mux10(\MEMTOREG|Mux10~1_combout ),
	.temp_iMemLoad_5(\EXMEM|temp_iMemLoad [5]),
	.alu_a_mux_output_21(\ALUAMUX|alu_a_mux_output[21]~64_combout ),
	.alu_a_mux_output_32(\ALUAMUX|alu_a_mux_output[3]~65_combout ),
	.always03(\FORWADUNIT|always0~19_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

mem_to_reg_mux MEMTOREG(
	.temp_dMemLoad_1(\MEMWB|temp_dMemLoad [1]),
	.temp_aluResult_1(\MEMWB|temp_aluResult [1]),
	.temp_memtoreg_0(\MEMWB|temp_memtoreg [0]),
	.temp_memtoreg_1(\MEMWB|temp_memtoreg [1]),
	.temp_npc_1(\MEMWB|temp_npc [1]),
	.Mux30(\MEMTOREG|Mux30~1_combout ),
	.temp_dMemLoad_0(\MEMWB|temp_dMemLoad [0]),
	.temp_aluResult_0(\MEMWB|temp_aluResult [0]),
	.temp_npc_0(\MEMWB|temp_npc [0]),
	.Mux31(\MEMTOREG|Mux31~1_combout ),
	.temp_dMemLoad_2(\MEMWB|temp_dMemLoad [2]),
	.temp_aluResult_2(\MEMWB|temp_aluResult [2]),
	.temp_npc_2(\MEMWB|temp_npc [2]),
	.Mux29(\MEMTOREG|Mux29~1_combout ),
	.temp_dMemLoad_4(\MEMWB|temp_dMemLoad [4]),
	.temp_aluResult_4(\MEMWB|temp_aluResult [4]),
	.temp_npc_4(\MEMWB|temp_npc [4]),
	.Mux27(\MEMTOREG|Mux27~1_combout ),
	.temp_dMemLoad_3(\MEMWB|temp_dMemLoad [3]),
	.temp_aluResult_3(\MEMWB|temp_aluResult [3]),
	.temp_npc_3(\MEMWB|temp_npc [3]),
	.Mux28(\MEMTOREG|Mux28~1_combout ),
	.temp_dMemLoad_8(\MEMWB|temp_dMemLoad [8]),
	.temp_aluResult_8(\MEMWB|temp_aluResult [8]),
	.temp_npc_8(\MEMWB|temp_npc [8]),
	.Mux23(\MEMTOREG|Mux23~1_combout ),
	.temp_dMemLoad_7(\MEMWB|temp_dMemLoad [7]),
	.temp_aluResult_7(\MEMWB|temp_aluResult [7]),
	.temp_npc_7(\MEMWB|temp_npc [7]),
	.Mux24(\MEMTOREG|Mux24~1_combout ),
	.temp_dMemLoad_6(\MEMWB|temp_dMemLoad [6]),
	.temp_aluResult_6(\MEMWB|temp_aluResult [6]),
	.temp_npc_6(\MEMWB|temp_npc [6]),
	.Mux25(\MEMTOREG|Mux25~1_combout ),
	.temp_dMemLoad_5(\MEMWB|temp_dMemLoad [5]),
	.temp_aluResult_5(\MEMWB|temp_aluResult [5]),
	.temp_npc_5(\MEMWB|temp_npc [5]),
	.Mux26(\MEMTOREG|Mux26~1_combout ),
	.temp_dMemLoad_16(\MEMWB|temp_dMemLoad [16]),
	.temp_upper16_16(\MEMWB|temp_upper16 [16]),
	.temp_aluResult_16(\MEMWB|temp_aluResult [16]),
	.temp_npc_16(\MEMWB|temp_npc [16]),
	.Mux15(\MEMTOREG|Mux15~1_combout ),
	.temp_dMemLoad_14(\MEMWB|temp_dMemLoad [14]),
	.temp_aluResult_14(\MEMWB|temp_aluResult [14]),
	.temp_npc_14(\MEMWB|temp_npc [14]),
	.Mux17(\MEMTOREG|Mux17~1_combout ),
	.temp_dMemLoad_15(\MEMWB|temp_dMemLoad [15]),
	.temp_aluResult_15(\MEMWB|temp_aluResult [15]),
	.temp_npc_15(\MEMWB|temp_npc [15]),
	.Mux16(\MEMTOREG|Mux16~1_combout ),
	.temp_dMemLoad_13(\MEMWB|temp_dMemLoad [13]),
	.temp_aluResult_13(\MEMWB|temp_aluResult [13]),
	.temp_npc_13(\MEMWB|temp_npc [13]),
	.Mux18(\MEMTOREG|Mux18~1_combout ),
	.temp_dMemLoad_12(\MEMWB|temp_dMemLoad [12]),
	.temp_aluResult_12(\MEMWB|temp_aluResult [12]),
	.temp_npc_12(\MEMWB|temp_npc [12]),
	.Mux19(\MEMTOREG|Mux19~1_combout ),
	.temp_dMemLoad_10(\MEMWB|temp_dMemLoad [10]),
	.temp_aluResult_10(\MEMWB|temp_aluResult [10]),
	.temp_npc_10(\MEMWB|temp_npc [10]),
	.Mux21(\MEMTOREG|Mux21~1_combout ),
	.temp_dMemLoad_11(\MEMWB|temp_dMemLoad [11]),
	.temp_aluResult_11(\MEMWB|temp_aluResult [11]),
	.temp_npc_11(\MEMWB|temp_npc [11]),
	.Mux20(\MEMTOREG|Mux20~1_combout ),
	.temp_dMemLoad_9(\MEMWB|temp_dMemLoad [9]),
	.temp_aluResult_9(\MEMWB|temp_aluResult [9]),
	.temp_npc_9(\MEMWB|temp_npc [9]),
	.Mux22(\MEMTOREG|Mux22~1_combout ),
	.temp_upper16_31(\MEMWB|temp_upper16 [31]),
	.temp_dMemLoad_31(\MEMWB|temp_dMemLoad [31]),
	.temp_aluResult_31(\MEMWB|temp_aluResult [31]),
	.temp_npc_31(\MEMWB|temp_npc [31]),
	.Mux0(\MEMTOREG|Mux0~1_combout ),
	.temp_dMemLoad_30(\MEMWB|temp_dMemLoad [30]),
	.temp_upper16_30(\MEMWB|temp_upper16 [30]),
	.temp_aluResult_30(\MEMWB|temp_aluResult [30]),
	.temp_npc_30(\MEMWB|temp_npc [30]),
	.Mux1(\MEMTOREG|Mux1~1_combout ),
	.temp_upper16_29(\MEMWB|temp_upper16 [29]),
	.temp_dMemLoad_29(\MEMWB|temp_dMemLoad [29]),
	.temp_aluResult_29(\MEMWB|temp_aluResult [29]),
	.temp_npc_29(\MEMWB|temp_npc [29]),
	.Mux2(\MEMTOREG|Mux2~1_combout ),
	.temp_upper16_26(\MEMWB|temp_upper16 [26]),
	.temp_dMemLoad_26(\MEMWB|temp_dMemLoad [26]),
	.temp_aluResult_26(\MEMWB|temp_aluResult [26]),
	.temp_npc_26(\MEMWB|temp_npc [26]),
	.Mux5(\MEMTOREG|Mux5~1_combout ),
	.temp_dMemLoad_25(\MEMWB|temp_dMemLoad [25]),
	.temp_upper16_25(\MEMWB|temp_upper16 [25]),
	.temp_aluResult_25(\MEMWB|temp_aluResult [25]),
	.temp_npc_25(\MEMWB|temp_npc [25]),
	.Mux6(\MEMTOREG|Mux6~1_combout ),
	.temp_dMemLoad_28(\MEMWB|temp_dMemLoad [28]),
	.temp_upper16_28(\MEMWB|temp_upper16 [28]),
	.temp_aluResult_28(\MEMWB|temp_aluResult [28]),
	.temp_npc_28(\MEMWB|temp_npc [28]),
	.Mux3(\MEMTOREG|Mux3~1_combout ),
	.temp_upper16_27(\MEMWB|temp_upper16 [27]),
	.temp_dMemLoad_27(\MEMWB|temp_dMemLoad [27]),
	.temp_aluResult_27(\MEMWB|temp_aluResult [27]),
	.temp_npc_27(\MEMWB|temp_npc [27]),
	.Mux4(\MEMTOREG|Mux4~1_combout ),
	.temp_upper16_17(\MEMWB|temp_upper16 [17]),
	.temp_dMemLoad_17(\MEMWB|temp_dMemLoad [17]),
	.temp_aluResult_17(\MEMWB|temp_aluResult [17]),
	.temp_npc_17(\MEMWB|temp_npc [17]),
	.Mux14(\MEMTOREG|Mux14~1_combout ),
	.temp_upper16_20(\MEMWB|temp_upper16 [20]),
	.temp_dMemLoad_20(\MEMWB|temp_dMemLoad [20]),
	.temp_aluResult_20(\MEMWB|temp_aluResult [20]),
	.temp_npc_20(\MEMWB|temp_npc [20]),
	.Mux11(\MEMTOREG|Mux11~1_combout ),
	.temp_dMemLoad_19(\MEMWB|temp_dMemLoad [19]),
	.temp_upper16_19(\MEMWB|temp_upper16 [19]),
	.temp_aluResult_19(\MEMWB|temp_aluResult [19]),
	.temp_npc_19(\MEMWB|temp_npc [19]),
	.Mux12(\MEMTOREG|Mux12~1_combout ),
	.temp_dMemLoad_18(\MEMWB|temp_dMemLoad [18]),
	.temp_upper16_18(\MEMWB|temp_upper16 [18]),
	.temp_aluResult_18(\MEMWB|temp_aluResult [18]),
	.temp_npc_18(\MEMWB|temp_npc [18]),
	.Mux13(\MEMTOREG|Mux13~1_combout ),
	.temp_upper16_24(\MEMWB|temp_upper16 [24]),
	.temp_dMemLoad_24(\MEMWB|temp_dMemLoad [24]),
	.temp_aluResult_24(\MEMWB|temp_aluResult [24]),
	.temp_npc_24(\MEMWB|temp_npc [24]),
	.Mux7(\MEMTOREG|Mux7~1_combout ),
	.temp_dMemLoad_23(\MEMWB|temp_dMemLoad [23]),
	.temp_upper16_23(\MEMWB|temp_upper16 [23]),
	.temp_aluResult_23(\MEMWB|temp_aluResult [23]),
	.temp_npc_23(\MEMWB|temp_npc [23]),
	.Mux8(\MEMTOREG|Mux8~1_combout ),
	.temp_upper16_22(\MEMWB|temp_upper16 [22]),
	.temp_dMemLoad_22(\MEMWB|temp_dMemLoad [22]),
	.temp_aluResult_22(\MEMWB|temp_aluResult [22]),
	.temp_npc_22(\MEMWB|temp_npc [22]),
	.Mux9(\MEMTOREG|Mux9~1_combout ),
	.temp_dMemLoad_21(\MEMWB|temp_dMemLoad [21]),
	.temp_upper16_21(\MEMWB|temp_upper16 [21]),
	.temp_aluResult_21(\MEMWB|temp_aluResult [21]),
	.temp_npc_21(\MEMWB|temp_npc [21]),
	.Mux10(\MEMTOREG|Mux10~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

alu_source_mux alusourceMUX(
	.temp_signzerovalue_output_16(\IDEX|temp_signzerovalue_output [16]),
	.temp_imemload_output_1(\IDEX|temp_imemload_output [1]),
	.temp_imemload_output_7(\IDEX|temp_imemload_output [7]),
	.temp_ALUsrc_output_1(\IDEX|temp_ALUsrc_output [1]),
	.temp_ALUsrc_output_0(\IDEX|temp_ALUsrc_output [0]),
	.Mux30(\alusourceMUX|Mux30~0_combout ),
	.alu_b_mux_output_1(\ALUBMUX|alu_b_mux_output[1]~0_combout ),
	.alu_b_mux_output_11(\ALUBMUX|alu_b_mux_output[1]~1_combout ),
	.Mux16(\alusourceMUX|Mux16~0_combout ),
	.Mux301(\alusourceMUX|Mux30~1_combout ),
	.alu_b_mux_output_0(\ALUBMUX|alu_b_mux_output[0]~2_combout ),
	.temp_imemload_output_0(\IDEX|temp_imemload_output [0]),
	.temp_imemload_output_6(\IDEX|temp_imemload_output [6]),
	.Mux31(\alusourceMUX|Mux31~0_combout ),
	.alu_b_mux_output_01(\ALUBMUX|alu_b_mux_output[0]~3_combout ),
	.Mux311(\alusourceMUX|Mux31~1_combout ),
	.temp_imemload_output_2(\IDEX|temp_imemload_output [2]),
	.temp_imemload_output_8(\IDEX|temp_imemload_output [8]),
	.Mux29(\alusourceMUX|Mux29~0_combout ),
	.alu_b_mux_output_2(\ALUBMUX|alu_b_mux_output[2]~5_combout ),
	.Mux291(\alusourceMUX|Mux29~1_combout ),
	.temp_imemload_output_3(\IDEX|temp_imemload_output [3]),
	.temp_imemload_output_9(\IDEX|temp_imemload_output [9]),
	.Mux28(\alusourceMUX|Mux28~0_combout ),
	.alu_b_mux_output_3(\ALUBMUX|alu_b_mux_output[3]~7_combout ),
	.Mux281(\alusourceMUX|Mux28~1_combout ),
	.temp_imemload_output_4(\IDEX|temp_imemload_output [4]),
	.temp_imemload_output_10(\IDEX|temp_imemload_output [10]),
	.Mux27(\alusourceMUX|Mux27~0_combout ),
	.alu_b_mux_output_4(\ALUBMUX|alu_b_mux_output[4]~9_combout ),
	.Mux271(\alusourceMUX|Mux27~1_combout ),
	.alu_b_mux_output_15(\ALUBMUX|alu_b_mux_output[15]~11_combout ),
	.temp_imemload_output_15(\IDEX|temp_imemload_output [15]),
	.Mux161(\alusourceMUX|Mux16~1_combout ),
	.alu_b_mux_output_12(\ALUBMUX|alu_b_mux_output[12]~13_combout ),
	.temp_imemload_output_12(\IDEX|temp_imemload_output [12]),
	.Mux19(\alusourceMUX|Mux19~0_combout ),
	.alu_b_mux_output_27(\ALUBMUX|alu_b_mux_output[27]~16_combout ),
	.Mux4(\alusourceMUX|Mux4~0_combout ),
	.alu_b_mux_output_18(\ALUBMUX|alu_b_mux_output[18]~18_combout ),
	.Mux13(\alusourceMUX|Mux13~0_combout ),
	.alu_b_mux_output_17(\ALUBMUX|alu_b_mux_output[17]~20_combout ),
	.Mux14(\alusourceMUX|Mux14~0_combout ),
	.alu_b_mux_output_16(\ALUBMUX|alu_b_mux_output[16]~22_combout ),
	.Mux15(\alusourceMUX|Mux15~0_combout ),
	.alu_b_mux_output_31(\ALUBMUX|alu_b_mux_output[31]~24_combout ),
	.Mux0(\alusourceMUX|Mux0~0_combout ),
	.alu_b_mux_output_30(\ALUBMUX|alu_b_mux_output[30]~26_combout ),
	.Mux1(\alusourceMUX|Mux1~0_combout ),
	.alu_b_mux_output_29(\ALUBMUX|alu_b_mux_output[29]~28_combout ),
	.Mux2(\alusourceMUX|Mux2~0_combout ),
	.alu_b_mux_output_28(\ALUBMUX|alu_b_mux_output[28]~30_combout ),
	.Mux3(\alusourceMUX|Mux3~0_combout ),
	.alu_b_mux_output_26(\ALUBMUX|alu_b_mux_output[26]~32_combout ),
	.Mux5(\alusourceMUX|Mux5~0_combout ),
	.alu_b_mux_output_25(\ALUBMUX|alu_b_mux_output[25]~34_combout ),
	.Mux6(\alusourceMUX|Mux6~0_combout ),
	.alu_b_mux_output_24(\ALUBMUX|alu_b_mux_output[24]~36_combout ),
	.Mux7(\alusourceMUX|Mux7~0_combout ),
	.alu_b_mux_output_23(\ALUBMUX|alu_b_mux_output[23]~38_combout ),
	.Mux8(\alusourceMUX|Mux8~0_combout ),
	.alu_b_mux_output_22(\ALUBMUX|alu_b_mux_output[22]~40_combout ),
	.Mux9(\alusourceMUX|Mux9~0_combout ),
	.alu_b_mux_output_21(\ALUBMUX|alu_b_mux_output[21]~42_combout ),
	.Mux10(\alusourceMUX|Mux10~0_combout ),
	.alu_b_mux_output_20(\ALUBMUX|alu_b_mux_output[20]~44_combout ),
	.Mux11(\alusourceMUX|Mux11~0_combout ),
	.alu_b_mux_output_19(\ALUBMUX|alu_b_mux_output[19]~46_combout ),
	.Mux12(\alusourceMUX|Mux12~0_combout ),
	.temp_imemload_output_14(\IDEX|temp_imemload_output [14]),
	.Mux17(\alusourceMUX|Mux17~0_combout ),
	.alu_b_mux_output_10(\ALUBMUX|alu_b_mux_output[10]~48_combout ),
	.Mux21(\alusourceMUX|Mux21~0_combout ),
	.alu_b_mux_output_14(\ALUBMUX|alu_b_mux_output[14]~50_combout ),
	.alu_b_mux_output_9(\ALUBMUX|alu_b_mux_output[9]~52_combout ),
	.Mux22(\alusourceMUX|Mux22~0_combout ),
	.alu_b_mux_output_8(\ALUBMUX|alu_b_mux_output[8]~54_combout ),
	.Mux23(\alusourceMUX|Mux23~0_combout ),
	.alu_b_mux_output_7(\ALUBMUX|alu_b_mux_output[7]~56_combout ),
	.Mux24(\alusourceMUX|Mux24~0_combout ),
	.alu_b_mux_output_6(\ALUBMUX|alu_b_mux_output[6]~58_combout ),
	.Mux25(\alusourceMUX|Mux25~0_combout ),
	.alu_b_mux_output_5(\ALUBMUX|alu_b_mux_output[5]~60_combout ),
	.temp_imemload_output_5(\IDEX|temp_imemload_output [5]),
	.Mux26(\alusourceMUX|Mux26~0_combout ),
	.alu_b_mux_output_13(\ALUBMUX|alu_b_mux_output[13]~62_combout ),
	.temp_imemload_output_13(\IDEX|temp_imemload_output [13]),
	.Mux18(\alusourceMUX|Mux18~0_combout ),
	.alu_b_mux_output_111(\ALUBMUX|alu_b_mux_output[11]~64_combout ),
	.temp_imemload_output_11(\IDEX|temp_imemload_output [11]),
	.Mux20(\alusourceMUX|Mux20~0_combout ),
	.Mux171(\alusourceMUX|Mux17~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

extender EXTENDER(
	.temp_imemload_output_31(\IFID|temp_imemload_output [31]),
	.temp_imemload_output_30(\IFID|temp_imemload_output [30]),
	.Equal3(\CONTROLUNIT|Equal3~0_combout ),
	.temp_branch_output(\IDEX|temp_branch_output~0_combout ),
	.temp_imemload_output_15(\IFID|temp_imemload_output [15]),
	.Equal31(\CONTROLUNIT|Equal3~9_combout ),
	.extended_imm_16(\EXTENDER|extended_imm[16]~0_combout ),
	.temp_ALUsrc_output(\IDEX|temp_ALUsrc_output~3_combout ),
	.WideOr5(\CONTROLUNIT|WideOr5~0_combout ),
	.extended_imm_161(\EXTENDER|extended_imm[16]~2_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

npc_mux NPCMUX(
	.temp_zeroFlag(\EXMEM|temp_zeroFlag~q ),
	.branch_count_output_2(\branch_count_output[2]~0_combout ),
	.pc_count_four_output_2(\pc_count_four_output[2]~0_combout ),
	.pc_count_four_output_3(\pc_count_four_output[3]~2_combout ),
	.branch_count_output_3(\branch_count_output[3]~2_combout ),
	.pc_count_four_output_4(\pc_count_four_output[4]~4_combout ),
	.pc_count_four_output_5(\pc_count_four_output[5]~6_combout ),
	.branch_count_output_4(\branch_count_output[4]~4_combout ),
	.branch_count_output_5(\branch_count_output[5]~6_combout ),
	.pc_count_four_output_6(\pc_count_four_output[6]~8_combout ),
	.pc_count_four_output_7(\pc_count_four_output[7]~10_combout ),
	.branch_count_output_6(\branch_count_output[6]~8_combout ),
	.branch_count_output_7(\branch_count_output[7]~10_combout ),
	.pc_count_four_output_8(\pc_count_four_output[8]~12_combout ),
	.pc_count_four_output_9(\pc_count_four_output[9]~14_combout ),
	.branch_count_output_8(\branch_count_output[8]~12_combout ),
	.branch_count_output_9(\branch_count_output[9]~14_combout ),
	.pc_count_four_output_10(\pc_count_four_output[10]~16_combout ),
	.pc_count_four_output_11(\pc_count_four_output[11]~18_combout ),
	.branch_count_output_10(\branch_count_output[10]~16_combout ),
	.branch_count_output_11(\branch_count_output[11]~18_combout ),
	.pc_count_four_output_12(\pc_count_four_output[12]~20_combout ),
	.pc_count_four_output_13(\pc_count_four_output[13]~22_combout ),
	.branch_count_output_12(\branch_count_output[12]~20_combout ),
	.branch_count_output_13(\branch_count_output[13]~22_combout ),
	.pc_count_four_output_14(\pc_count_four_output[14]~24_combout ),
	.pc_count_four_output_15(\pc_count_four_output[15]~26_combout ),
	.branch_count_output_14(\branch_count_output[14]~24_combout ),
	.branch_count_output_15(\branch_count_output[15]~26_combout ),
	.pc_count_four_output_16(\pc_count_four_output[16]~28_combout ),
	.pc_count_four_output_17(\pc_count_four_output[17]~30_combout ),
	.branch_count_output_16(\branch_count_output[16]~28_combout ),
	.branch_count_output_17(\branch_count_output[17]~30_combout ),
	.pc_count_four_output_18(\pc_count_four_output[18]~32_combout ),
	.pc_count_four_output_19(\pc_count_four_output[19]~34_combout ),
	.branch_count_output_18(\branch_count_output[18]~32_combout ),
	.branch_count_output_19(\branch_count_output[19]~34_combout ),
	.branch_count_output_20(\branch_count_output[20]~36_combout ),
	.pc_count_four_output_20(\pc_count_four_output[20]~36_combout ),
	.pc_count_four_output_21(\pc_count_four_output[21]~38_combout ),
	.branch_count_output_21(\branch_count_output[21]~38_combout ),
	.pc_count_four_output_22(\pc_count_four_output[22]~40_combout ),
	.pc_count_four_output_23(\pc_count_four_output[23]~42_combout ),
	.branch_count_output_22(\branch_count_output[22]~40_combout ),
	.branch_count_output_23(\branch_count_output[23]~42_combout ),
	.pc_count_four_output_24(\pc_count_four_output[24]~44_combout ),
	.pc_count_four_output_25(\pc_count_four_output[25]~46_combout ),
	.branch_count_output_24(\branch_count_output[24]~44_combout ),
	.branch_count_output_25(\branch_count_output[25]~46_combout ),
	.branch_count_output_26(\branch_count_output[26]~48_combout ),
	.pc_count_four_output_26(\pc_count_four_output[26]~48_combout ),
	.pc_count_four_output_27(\pc_count_four_output[27]~50_combout ),
	.pc_count_four_output_28(\pc_count_four_output[28]~52_combout ),
	.branch_count_output_27(\branch_count_output[27]~50_combout ),
	.pc_count_four_output_29(\pc_count_four_output[29]~54_combout ),
	.branch_count_output_28(\branch_count_output[28]~52_combout ),
	.branch_count_output_29(\branch_count_output[29]~54_combout ),
	.pc_count_four_output_30(\pc_count_four_output[30]~56_combout ),
	.pc_count_four_output_31(\pc_count_four_output[31]~58_combout ),
	.branch_count_output_30(\branch_count_output[30]~56_combout ),
	.branch_count_output_31(\branch_count_output[31]~58_combout ),
	.pccount_1(pccount_1),
	.pccount_0(pccount_0),
	.temp_iMemLoad_0(\EXMEM|temp_iMemLoad [0]),
	.temp_iMemLoad_15(\EXMEM|temp_iMemLoad [15]),
	.temp_iMemLoad_14(\EXMEM|temp_iMemLoad [14]),
	.temp_iMemLoad_13(\EXMEM|temp_iMemLoad [13]),
	.temp_iMemLoad_10(\EXMEM|temp_iMemLoad [10]),
	.temp_iMemLoad_9(\EXMEM|temp_iMemLoad [9]),
	.temp_iMemLoad_12(\EXMEM|temp_iMemLoad [12]),
	.temp_iMemLoad_11(\EXMEM|temp_iMemLoad [11]),
	.temp_iMemLoad_1(\EXMEM|temp_iMemLoad [1]),
	.temp_iMemLoad_4(\EXMEM|temp_iMemLoad [4]),
	.temp_iMemLoad_3(\EXMEM|temp_iMemLoad [3]),
	.temp_iMemLoad_2(\EXMEM|temp_iMemLoad [2]),
	.temp_iMemLoad_8(\EXMEM|temp_iMemLoad [8]),
	.temp_iMemLoad_7(\EXMEM|temp_iMemLoad [7]),
	.temp_iMemLoad_6(\EXMEM|temp_iMemLoad [6]),
	.temp_iMemLoad_5(\EXMEM|temp_iMemLoad [5]),
	.temp_branchSelect(\EXMEM|temp_branchSelect~q ),
	.temp_rdat1_1(\EXMEM|temp_rdat1 [1]),
	.temp_npc_1(\EXMEM|temp_npc [1]),
	.temp_pcselect_1(\EXMEM|temp_pcselect [1]),
	.temp_pcselect_0(\EXMEM|temp_pcselect [0]),
	.Mux30(\NPCMUX|Mux30~1_combout ),
	.temp_rdat1_0(\EXMEM|temp_rdat1 [0]),
	.temp_npc_0(\EXMEM|temp_npc [0]),
	.Mux31(\NPCMUX|Mux31~2_combout ),
	.temp_rdat1_2(\EXMEM|temp_rdat1 [2]),
	.Mux29(\NPCMUX|Mux29~1_combout ),
	.temp_rdat1_3(\EXMEM|temp_rdat1 [3]),
	.Mux28(\NPCMUX|Mux28~1_combout ),
	.temp_rdat1_5(\EXMEM|temp_rdat1 [5]),
	.Mux26(\NPCMUX|Mux26~1_combout ),
	.temp_rdat1_4(\EXMEM|temp_rdat1 [4]),
	.Mux27(\NPCMUX|Mux27~1_combout ),
	.temp_rdat1_7(\EXMEM|temp_rdat1 [7]),
	.Mux24(\NPCMUX|Mux24~1_combout ),
	.temp_rdat1_6(\EXMEM|temp_rdat1 [6]),
	.Mux25(\NPCMUX|Mux25~1_combout ),
	.temp_rdat1_9(\EXMEM|temp_rdat1 [9]),
	.Mux22(\NPCMUX|Mux22~1_combout ),
	.temp_rdat1_8(\EXMEM|temp_rdat1 [8]),
	.Mux23(\NPCMUX|Mux23~1_combout ),
	.temp_rdat1_11(\EXMEM|temp_rdat1 [11]),
	.Mux20(\NPCMUX|Mux20~1_combout ),
	.temp_rdat1_10(\EXMEM|temp_rdat1 [10]),
	.Mux21(\NPCMUX|Mux21~1_combout ),
	.temp_rdat1_13(\EXMEM|temp_rdat1 [13]),
	.Mux18(\NPCMUX|Mux18~1_combout ),
	.temp_rdat1_12(\EXMEM|temp_rdat1 [12]),
	.Mux19(\NPCMUX|Mux19~1_combout ),
	.temp_rdat1_15(\EXMEM|temp_rdat1 [15]),
	.Mux16(\NPCMUX|Mux16~1_combout ),
	.temp_rdat1_14(\EXMEM|temp_rdat1 [14]),
	.Mux17(\NPCMUX|Mux17~1_combout ),
	.temp_rdat1_17(\EXMEM|temp_rdat1 [17]),
	.Mux14(\NPCMUX|Mux14~1_combout ),
	.temp_rdat1_16(\EXMEM|temp_rdat1 [16]),
	.Mux15(\NPCMUX|Mux15~1_combout ),
	.temp_rdat1_19(\EXMEM|temp_rdat1 [19]),
	.temp_iMemLoad_17(\EXMEM|temp_iMemLoad [17]),
	.Mux12(\NPCMUX|Mux12~1_combout ),
	.temp_rdat1_18(\EXMEM|temp_rdat1 [18]),
	.temp_iMemLoad_16(\EXMEM|temp_iMemLoad [16]),
	.Mux13(\NPCMUX|Mux13~1_combout ),
	.temp_rdat1_20(\EXMEM|temp_rdat1 [20]),
	.temp_iMemLoad_18(\EXMEM|temp_iMemLoad [18]),
	.Mux11(\NPCMUX|Mux11~1_combout ),
	.temp_rdat1_21(\EXMEM|temp_rdat1 [21]),
	.temp_iMemLoad_19(\EXMEM|temp_iMemLoad [19]),
	.Mux10(\NPCMUX|Mux10~1_combout ),
	.temp_rdat1_23(\EXMEM|temp_rdat1 [23]),
	.temp_iMemLoad_21(\EXMEM|temp_iMemLoad [21]),
	.Mux8(\NPCMUX|Mux8~1_combout ),
	.temp_rdat1_22(\EXMEM|temp_rdat1 [22]),
	.temp_iMemLoad_20(\EXMEM|temp_iMemLoad [20]),
	.Mux9(\NPCMUX|Mux9~1_combout ),
	.temp_rdat1_25(\EXMEM|temp_rdat1 [25]),
	.temp_iMemLoad_23(\EXMEM|temp_iMemLoad [23]),
	.Mux6(\NPCMUX|Mux6~1_combout ),
	.temp_rdat1_24(\EXMEM|temp_rdat1 [24]),
	.temp_iMemLoad_22(\EXMEM|temp_iMemLoad [22]),
	.Mux7(\NPCMUX|Mux7~1_combout ),
	.temp_rdat1_26(\EXMEM|temp_rdat1 [26]),
	.Mux5(\NPCMUX|Mux5~1_combout ),
	.temp_rdat1_27(\EXMEM|temp_rdat1 [27]),
	.Mux4(\NPCMUX|Mux4~1_combout ),
	.temp_rdat1_29(\EXMEM|temp_rdat1 [29]),
	.Mux2(\NPCMUX|Mux2~1_combout ),
	.temp_rdat1_28(\EXMEM|temp_rdat1 [28]),
	.Mux3(\NPCMUX|Mux3~3_combout ),
	.temp_rdat1_31(\EXMEM|temp_rdat1 [31]),
	.Mux0(\NPCMUX|Mux0~1_combout ),
	.temp_rdat1_30(\EXMEM|temp_rdat1 [30]),
	.Mux1(\NPCMUX|Mux1~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

mem_wb_latch MEMWB(
	.temp_branchDest_0(\EXMEM|temp_branchDest [0]),
	.temp_branchDest_4(\EXMEM|temp_branchDest [4]),
	.temp_branchDest_3(\EXMEM|temp_branchDest [3]),
	.temp_branchDest_2(\EXMEM|temp_branchDest [2]),
	.temp_branchDest_1(\EXMEM|temp_branchDest [1]),
	.temp_aluResult_1(temp_aluResult_1),
	.temp_aluResult_0(temp_aluResult_0),
	.temp_aluResult_2(temp_aluResult_2),
	.temp_aluResult_3(temp_aluResult_3),
	.temp_aluResult_5(temp_aluResult_5),
	.temp_aluResult_4(temp_aluResult_4),
	.temp_aluResult_7(temp_aluResult_7),
	.temp_aluResult_6(temp_aluResult_6),
	.temp_aluResult_9(temp_aluResult_9),
	.temp_aluResult_8(temp_aluResult_8),
	.temp_aluResult_11(temp_aluResult_11),
	.temp_aluResult_10(temp_aluResult_10),
	.temp_aluResult_13(temp_aluResult_13),
	.temp_aluResult_12(temp_aluResult_12),
	.temp_aluResult_15(temp_aluResult_15),
	.temp_aluResult_14(temp_aluResult_14),
	.temp_aluResult_17(temp_aluResult_17),
	.temp_aluResult_16(temp_aluResult_16),
	.temp_aluResult_19(temp_aluResult_19),
	.temp_aluResult_18(temp_aluResult_18),
	.temp_aluResult_20(temp_aluResult_20),
	.temp_aluResult_21(temp_aluResult_21),
	.temp_aluResult_23(temp_aluResult_23),
	.temp_aluResult_22(temp_aluResult_22),
	.temp_aluResult_25(temp_aluResult_25),
	.temp_aluResult_24(temp_aluResult_24),
	.temp_aluResult_26(temp_aluResult_26),
	.temp_aluResult_27(temp_aluResult_27),
	.temp_aluResult_29(temp_aluResult_29),
	.temp_aluResult_28(temp_aluResult_28),
	.temp_aluResult_31(temp_aluResult_31),
	.temp_aluResult_30(temp_aluResult_30),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.temp_regwrite1(\EXMEM|temp_regwrite~q ),
	.temp_memtoreg_0(\EXMEM|temp_memtoreg [0]),
	.temp_memtoreg_1(\EXMEM|temp_memtoreg [1]),
	.temp_regwrite2(\MEMWB|temp_regwrite~q ),
	.temp_branchDest_11(\MEMWB|temp_branchDest [1]),
	.temp_branchDest_01(\MEMWB|temp_branchDest [0]),
	.temp_branchDest_31(\MEMWB|temp_branchDest [3]),
	.temp_branchDest_21(\MEMWB|temp_branchDest [2]),
	.temp_branchDest_41(\MEMWB|temp_branchDest [4]),
	.temp_dMemLoad_1(\MEMWB|temp_dMemLoad [1]),
	.temp_aluResult_110(\MEMWB|temp_aluResult [1]),
	.temp_memtoreg_01(\MEMWB|temp_memtoreg [0]),
	.temp_memtoreg_11(\MEMWB|temp_memtoreg [1]),
	.temp_npc_1(\MEMWB|temp_npc [1]),
	.temp_dMemLoad_0(\MEMWB|temp_dMemLoad [0]),
	.temp_aluResult_01(\MEMWB|temp_aluResult [0]),
	.temp_npc_0(\MEMWB|temp_npc [0]),
	.temp_dMemLoad_2(\MEMWB|temp_dMemLoad [2]),
	.temp_aluResult_210(\MEMWB|temp_aluResult [2]),
	.temp_npc_2(\MEMWB|temp_npc [2]),
	.temp_dMemLoad_4(\MEMWB|temp_dMemLoad [4]),
	.temp_aluResult_41(\MEMWB|temp_aluResult [4]),
	.temp_npc_4(\MEMWB|temp_npc [4]),
	.temp_dMemLoad_3(\MEMWB|temp_dMemLoad [3]),
	.temp_aluResult_32(\MEMWB|temp_aluResult [3]),
	.temp_npc_3(\MEMWB|temp_npc [3]),
	.temp_dMemLoad_8(\MEMWB|temp_dMemLoad [8]),
	.temp_aluResult_81(\MEMWB|temp_aluResult [8]),
	.temp_npc_8(\MEMWB|temp_npc [8]),
	.temp_dMemLoad_7(\MEMWB|temp_dMemLoad [7]),
	.temp_aluResult_71(\MEMWB|temp_aluResult [7]),
	.temp_npc_7(\MEMWB|temp_npc [7]),
	.temp_dMemLoad_6(\MEMWB|temp_dMemLoad [6]),
	.temp_aluResult_61(\MEMWB|temp_aluResult [6]),
	.temp_npc_6(\MEMWB|temp_npc [6]),
	.temp_dMemLoad_5(\MEMWB|temp_dMemLoad [5]),
	.temp_aluResult_51(\MEMWB|temp_aluResult [5]),
	.temp_npc_5(\MEMWB|temp_npc [5]),
	.temp_dMemLoad_16(\MEMWB|temp_dMemLoad [16]),
	.temp_upper16_16(\MEMWB|temp_upper16 [16]),
	.temp_aluResult_161(\MEMWB|temp_aluResult [16]),
	.temp_npc_16(\MEMWB|temp_npc [16]),
	.temp_iMemLoad_0(\EXMEM|temp_iMemLoad [0]),
	.temp_dMemLoad_14(\MEMWB|temp_dMemLoad [14]),
	.temp_aluResult_141(\MEMWB|temp_aluResult [14]),
	.temp_npc_14(\MEMWB|temp_npc [14]),
	.temp_dMemLoad_15(\MEMWB|temp_dMemLoad [15]),
	.temp_aluResult_151(\MEMWB|temp_aluResult [15]),
	.temp_npc_15(\MEMWB|temp_npc [15]),
	.temp_dMemLoad_13(\MEMWB|temp_dMemLoad [13]),
	.temp_aluResult_131(\MEMWB|temp_aluResult [13]),
	.temp_npc_13(\MEMWB|temp_npc [13]),
	.temp_dMemLoad_12(\MEMWB|temp_dMemLoad [12]),
	.temp_aluResult_121(\MEMWB|temp_aluResult [12]),
	.temp_npc_12(\MEMWB|temp_npc [12]),
	.temp_dMemLoad_10(\MEMWB|temp_dMemLoad [10]),
	.temp_aluResult_101(\MEMWB|temp_aluResult [10]),
	.temp_npc_10(\MEMWB|temp_npc [10]),
	.temp_dMemLoad_11(\MEMWB|temp_dMemLoad [11]),
	.temp_aluResult_111(\MEMWB|temp_aluResult [11]),
	.temp_npc_11(\MEMWB|temp_npc [11]),
	.temp_dMemLoad_9(\MEMWB|temp_dMemLoad [9]),
	.temp_aluResult_91(\MEMWB|temp_aluResult [9]),
	.temp_npc_9(\MEMWB|temp_npc [9]),
	.temp_upper16_31(\MEMWB|temp_upper16 [31]),
	.temp_dMemLoad_31(\MEMWB|temp_dMemLoad [31]),
	.temp_aluResult_311(\MEMWB|temp_aluResult [31]),
	.temp_npc_31(\MEMWB|temp_npc [31]),
	.temp_iMemLoad_15(\EXMEM|temp_iMemLoad [15]),
	.temp_dMemLoad_30(\MEMWB|temp_dMemLoad [30]),
	.temp_upper16_30(\MEMWB|temp_upper16 [30]),
	.temp_aluResult_301(\MEMWB|temp_aluResult [30]),
	.temp_npc_30(\MEMWB|temp_npc [30]),
	.temp_iMemLoad_14(\EXMEM|temp_iMemLoad [14]),
	.temp_upper16_29(\MEMWB|temp_upper16 [29]),
	.temp_dMemLoad_29(\MEMWB|temp_dMemLoad [29]),
	.temp_aluResult_291(\MEMWB|temp_aluResult [29]),
	.temp_npc_29(\MEMWB|temp_npc [29]),
	.temp_iMemLoad_13(\EXMEM|temp_iMemLoad [13]),
	.temp_upper16_26(\MEMWB|temp_upper16 [26]),
	.temp_dMemLoad_26(\MEMWB|temp_dMemLoad [26]),
	.temp_aluResult_261(\MEMWB|temp_aluResult [26]),
	.temp_npc_26(\MEMWB|temp_npc [26]),
	.temp_iMemLoad_10(\EXMEM|temp_iMemLoad [10]),
	.temp_dMemLoad_25(\MEMWB|temp_dMemLoad [25]),
	.temp_upper16_25(\MEMWB|temp_upper16 [25]),
	.temp_aluResult_251(\MEMWB|temp_aluResult [25]),
	.temp_npc_25(\MEMWB|temp_npc [25]),
	.temp_iMemLoad_9(\EXMEM|temp_iMemLoad [9]),
	.temp_dMemLoad_28(\MEMWB|temp_dMemLoad [28]),
	.temp_upper16_28(\MEMWB|temp_upper16 [28]),
	.temp_aluResult_281(\MEMWB|temp_aluResult [28]),
	.temp_npc_28(\MEMWB|temp_npc [28]),
	.temp_iMemLoad_12(\EXMEM|temp_iMemLoad [12]),
	.temp_upper16_27(\MEMWB|temp_upper16 [27]),
	.temp_dMemLoad_27(\MEMWB|temp_dMemLoad [27]),
	.temp_aluResult_271(\MEMWB|temp_aluResult [27]),
	.temp_npc_27(\MEMWB|temp_npc [27]),
	.temp_iMemLoad_11(\EXMEM|temp_iMemLoad [11]),
	.temp_upper16_17(\MEMWB|temp_upper16 [17]),
	.temp_dMemLoad_17(\MEMWB|temp_dMemLoad [17]),
	.temp_aluResult_171(\MEMWB|temp_aluResult [17]),
	.temp_npc_17(\MEMWB|temp_npc [17]),
	.temp_iMemLoad_1(\EXMEM|temp_iMemLoad [1]),
	.temp_upper16_20(\MEMWB|temp_upper16 [20]),
	.temp_dMemLoad_20(\MEMWB|temp_dMemLoad [20]),
	.temp_aluResult_201(\MEMWB|temp_aluResult [20]),
	.temp_npc_20(\MEMWB|temp_npc [20]),
	.temp_iMemLoad_4(\EXMEM|temp_iMemLoad [4]),
	.temp_dMemLoad_19(\MEMWB|temp_dMemLoad [19]),
	.temp_upper16_19(\MEMWB|temp_upper16 [19]),
	.temp_aluResult_191(\MEMWB|temp_aluResult [19]),
	.temp_npc_19(\MEMWB|temp_npc [19]),
	.temp_iMemLoad_3(\EXMEM|temp_iMemLoad [3]),
	.temp_dMemLoad_18(\MEMWB|temp_dMemLoad [18]),
	.temp_upper16_18(\MEMWB|temp_upper16 [18]),
	.temp_aluResult_181(\MEMWB|temp_aluResult [18]),
	.temp_npc_18(\MEMWB|temp_npc [18]),
	.temp_iMemLoad_2(\EXMEM|temp_iMemLoad [2]),
	.temp_upper16_24(\MEMWB|temp_upper16 [24]),
	.temp_dMemLoad_24(\MEMWB|temp_dMemLoad [24]),
	.temp_aluResult_241(\MEMWB|temp_aluResult [24]),
	.temp_npc_24(\MEMWB|temp_npc [24]),
	.temp_iMemLoad_8(\EXMEM|temp_iMemLoad [8]),
	.temp_dMemLoad_23(\MEMWB|temp_dMemLoad [23]),
	.temp_upper16_23(\MEMWB|temp_upper16 [23]),
	.temp_aluResult_231(\MEMWB|temp_aluResult [23]),
	.temp_npc_23(\MEMWB|temp_npc [23]),
	.temp_iMemLoad_7(\EXMEM|temp_iMemLoad [7]),
	.temp_upper16_22(\MEMWB|temp_upper16 [22]),
	.temp_dMemLoad_22(\MEMWB|temp_dMemLoad [22]),
	.temp_aluResult_221(\MEMWB|temp_aluResult [22]),
	.temp_npc_22(\MEMWB|temp_npc [22]),
	.temp_iMemLoad_6(\EXMEM|temp_iMemLoad [6]),
	.temp_dMemLoad_21(\MEMWB|temp_dMemLoad [21]),
	.temp_upper16_21(\MEMWB|temp_upper16 [21]),
	.temp_aluResult_211(\MEMWB|temp_aluResult [21]),
	.temp_npc_21(\MEMWB|temp_npc [21]),
	.temp_iMemLoad_5(\EXMEM|temp_iMemLoad [5]),
	.wen(\HAZARDUNIT|id_ex_wen~0_combout ),
	.temp_npc_110(\EXMEM|temp_npc [1]),
	.temp_npc_01(\EXMEM|temp_npc [0]),
	.temp_npc_210(\EXMEM|temp_npc [2]),
	.temp_npc_32(\EXMEM|temp_npc [3]),
	.temp_npc_51(\EXMEM|temp_npc [5]),
	.temp_npc_41(\EXMEM|temp_npc [4]),
	.temp_npc_71(\EXMEM|temp_npc [7]),
	.temp_npc_61(\EXMEM|temp_npc [6]),
	.temp_npc_91(\EXMEM|temp_npc [9]),
	.temp_npc_81(\EXMEM|temp_npc [8]),
	.temp_npc_111(\EXMEM|temp_npc [11]),
	.temp_npc_101(\EXMEM|temp_npc [10]),
	.temp_npc_131(\EXMEM|temp_npc [13]),
	.temp_npc_121(\EXMEM|temp_npc [12]),
	.temp_npc_151(\EXMEM|temp_npc [15]),
	.temp_npc_141(\EXMEM|temp_npc [14]),
	.temp_npc_171(\EXMEM|temp_npc [17]),
	.temp_npc_161(\EXMEM|temp_npc [16]),
	.temp_npc_191(\EXMEM|temp_npc [19]),
	.temp_npc_181(\EXMEM|temp_npc [18]),
	.temp_npc_201(\EXMEM|temp_npc [20]),
	.temp_npc_211(\EXMEM|temp_npc [21]),
	.temp_npc_231(\EXMEM|temp_npc [23]),
	.temp_npc_221(\EXMEM|temp_npc [22]),
	.temp_npc_251(\EXMEM|temp_npc [25]),
	.temp_npc_241(\EXMEM|temp_npc [24]),
	.temp_npc_261(\EXMEM|temp_npc [26]),
	.temp_npc_271(\EXMEM|temp_npc [27]),
	.temp_npc_291(\EXMEM|temp_npc [29]),
	.temp_npc_281(\EXMEM|temp_npc [28]),
	.temp_npc_311(\EXMEM|temp_npc [31]),
	.temp_npc_301(\EXMEM|temp_npc [30]),
	.CLK(CPUCLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

ex_mem_latch EXMEM(
	.temp_branchDest_0(\EXMEM|temp_branchDest [0]),
	.temp_branchDest_4(\EXMEM|temp_branchDest [4]),
	.temp_branchDest_3(\EXMEM|temp_branchDest [3]),
	.temp_branchDest_2(\EXMEM|temp_branchDest [2]),
	.temp_branchDest_1(\EXMEM|temp_branchDest [1]),
	.temp_signzerovalue_output_16(\IDEX|temp_signzerovalue_output [16]),
	.temp_zeroFlag1(\EXMEM|temp_zeroFlag~q ),
	.temp_halt_out_output(\IDEX|temp_halt_out_output~q ),
	.temp_aluResult_1(temp_aluResult_1),
	.temp_dmemWEN1(temp_dmemWEN),
	.temp_dmemREN1(temp_dmemREN),
	.temp_aluResult_0(temp_aluResult_0),
	.temp_aluResult_2(temp_aluResult_2),
	.temp_aluResult_3(temp_aluResult_3),
	.temp_aluResult_5(temp_aluResult_5),
	.temp_aluResult_4(temp_aluResult_4),
	.temp_aluResult_7(temp_aluResult_7),
	.temp_aluResult_6(temp_aluResult_6),
	.temp_aluResult_9(temp_aluResult_9),
	.temp_aluResult_8(temp_aluResult_8),
	.temp_aluResult_11(temp_aluResult_11),
	.temp_aluResult_10(temp_aluResult_10),
	.temp_aluResult_13(temp_aluResult_13),
	.temp_aluResult_12(temp_aluResult_12),
	.temp_aluResult_15(temp_aluResult_15),
	.temp_aluResult_14(temp_aluResult_14),
	.temp_aluResult_17(temp_aluResult_17),
	.temp_aluResult_16(temp_aluResult_16),
	.temp_aluResult_19(temp_aluResult_19),
	.temp_aluResult_18(temp_aluResult_18),
	.temp_aluResult_20(temp_aluResult_20),
	.temp_aluResult_21(temp_aluResult_21),
	.temp_aluResult_23(temp_aluResult_23),
	.temp_aluResult_22(temp_aluResult_22),
	.temp_aluResult_25(temp_aluResult_25),
	.temp_aluResult_24(temp_aluResult_24),
	.temp_aluResult_26(temp_aluResult_26),
	.temp_aluResult_27(temp_aluResult_27),
	.temp_aluResult_29(temp_aluResult_29),
	.temp_aluResult_28(temp_aluResult_28),
	.temp_aluResult_31(temp_aluResult_31),
	.temp_aluResult_30(temp_aluResult_30),
	.temp_halt_out1(\EXMEM|temp_halt_out~q ),
	.temp_rdat2_0(temp_rdat2_0),
	.temp_imemload_output_1(\IDEX|temp_imemload_output [1]),
	.temp_imemload_output_7(\IDEX|temp_imemload_output [7]),
	.temp_regwrite1(\EXMEM|temp_regwrite~q ),
	.temp_imemload_output_17(\IDEX|temp_imemload_output [17]),
	.temp_imemload_output_16(\IDEX|temp_imemload_output [16]),
	.temp_imemload_output_18(\IDEX|temp_imemload_output [18]),
	.temp_imemload_output_19(\IDEX|temp_imemload_output [19]),
	.temp_imemload_output_20(\IDEX|temp_imemload_output [20]),
	.temp_memtoreg_0(\EXMEM|temp_memtoreg [0]),
	.temp_memtoreg_1(\EXMEM|temp_memtoreg [1]),
	.alu_b_mux_output_1(\ALUBMUX|alu_b_mux_output[1]~0_combout ),
	.alu_b_mux_output_11(\ALUBMUX|alu_b_mux_output[1]~1_combout ),
	.temp_imemload_output_22(\IDEX|temp_imemload_output [22]),
	.temp_imemload_output_21(\IDEX|temp_imemload_output [21]),
	.temp_imemload_output_23(\IDEX|temp_imemload_output [23]),
	.alu_a_mux_output_1(\ALUAMUX|alu_a_mux_output[1]~1_combout ),
	.alu_b_mux_output_0(\ALUBMUX|alu_b_mux_output[0]~2_combout ),
	.temp_imemload_output_0(\IDEX|temp_imemload_output [0]),
	.temp_imemload_output_6(\IDEX|temp_imemload_output [6]),
	.alu_b_mux_output_01(\ALUBMUX|alu_b_mux_output[0]~3_combout ),
	.alu_a_mux_output_0(\ALUAMUX|alu_a_mux_output[0]~3_combout ),
	.alu_a_mux_output_2(\ALUAMUX|alu_a_mux_output[2]~5_combout ),
	.alu_a_mux_output_4(\ALUAMUX|alu_a_mux_output[4]~7_combout ),
	.alu_a_mux_output_3(\ALUAMUX|alu_a_mux_output[3]~8_combout ),
	.temp_imemload_output_2(\IDEX|temp_imemload_output [2]),
	.temp_imemload_output_8(\IDEX|temp_imemload_output [8]),
	.alu_b_mux_output_2(\ALUBMUX|alu_b_mux_output[2]~5_combout ),
	.alu_a_mux_output_8(\ALUAMUX|alu_a_mux_output[8]~11_combout ),
	.alu_a_mux_output_7(\ALUAMUX|alu_a_mux_output[7]~13_combout ),
	.alu_a_mux_output_6(\ALUAMUX|alu_a_mux_output[6]~15_combout ),
	.alu_a_mux_output_5(\ALUAMUX|alu_a_mux_output[5]~17_combout ),
	.temp_imemload_output_3(\IDEX|temp_imemload_output [3]),
	.temp_imemload_output_9(\IDEX|temp_imemload_output [9]),
	.alu_b_mux_output_3(\ALUBMUX|alu_b_mux_output[3]~7_combout ),
	.temp_iMemLoad_0(\EXMEM|temp_iMemLoad [0]),
	.alu_a_mux_output_16(\ALUAMUX|alu_a_mux_output[16]~20_combout ),
	.alu_a_mux_output_14(\ALUAMUX|alu_a_mux_output[14]~22_combout ),
	.alu_a_mux_output_15(\ALUAMUX|alu_a_mux_output[15]~24_combout ),
	.alu_a_mux_output_13(\ALUAMUX|alu_a_mux_output[13]~26_combout ),
	.alu_a_mux_output_12(\ALUAMUX|alu_a_mux_output[12]~28_combout ),
	.alu_a_mux_output_10(\ALUAMUX|alu_a_mux_output[10]~30_combout ),
	.alu_a_mux_output_11(\ALUAMUX|alu_a_mux_output[11]~32_combout ),
	.alu_a_mux_output_9(\ALUAMUX|alu_a_mux_output[9]~34_combout ),
	.temp_imemload_output_4(\IDEX|temp_imemload_output [4]),
	.temp_imemload_output_10(\IDEX|temp_imemload_output [10]),
	.alu_b_mux_output_4(\ALUBMUX|alu_b_mux_output[4]~9_combout ),
	.temp_iMemLoad_15(\EXMEM|temp_iMemLoad [15]),
	.alu_a_mux_output_31(\ALUAMUX|alu_a_mux_output[31]~36_combout ),
	.temp_iMemLoad_14(\EXMEM|temp_iMemLoad [14]),
	.alu_a_mux_output_30(\ALUAMUX|alu_a_mux_output[30]~38_combout ),
	.temp_iMemLoad_13(\EXMEM|temp_iMemLoad [13]),
	.alu_a_mux_output_29(\ALUAMUX|alu_a_mux_output[29]~40_combout ),
	.temp_iMemLoad_10(\EXMEM|temp_iMemLoad [10]),
	.alu_a_mux_output_26(\ALUAMUX|alu_a_mux_output[26]~42_combout ),
	.temp_iMemLoad_9(\EXMEM|temp_iMemLoad [9]),
	.alu_a_mux_output_25(\ALUAMUX|alu_a_mux_output[25]~44_combout ),
	.temp_iMemLoad_12(\EXMEM|temp_iMemLoad [12]),
	.alu_a_mux_output_28(\ALUAMUX|alu_a_mux_output[28]~46_combout ),
	.temp_iMemLoad_11(\EXMEM|temp_iMemLoad [11]),
	.alu_a_mux_output_27(\ALUAMUX|alu_a_mux_output[27]~48_combout ),
	.temp_iMemLoad_1(\EXMEM|temp_iMemLoad [1]),
	.alu_a_mux_output_17(\ALUAMUX|alu_a_mux_output[17]~50_combout ),
	.temp_iMemLoad_4(\EXMEM|temp_iMemLoad [4]),
	.alu_a_mux_output_20(\ALUAMUX|alu_a_mux_output[20]~52_combout ),
	.temp_iMemLoad_3(\EXMEM|temp_iMemLoad [3]),
	.alu_a_mux_output_19(\ALUAMUX|alu_a_mux_output[19]~54_combout ),
	.temp_iMemLoad_2(\EXMEM|temp_iMemLoad [2]),
	.alu_a_mux_output_18(\ALUAMUX|alu_a_mux_output[18]~56_combout ),
	.temp_iMemLoad_8(\EXMEM|temp_iMemLoad [8]),
	.alu_a_mux_output_24(\ALUAMUX|alu_a_mux_output[24]~58_combout ),
	.temp_iMemLoad_7(\EXMEM|temp_iMemLoad [7]),
	.alu_a_mux_output_23(\ALUAMUX|alu_a_mux_output[23]~60_combout ),
	.temp_iMemLoad_6(\EXMEM|temp_iMemLoad [6]),
	.alu_a_mux_output_22(\ALUAMUX|alu_a_mux_output[22]~62_combout ),
	.temp_iMemLoad_5(\EXMEM|temp_iMemLoad [5]),
	.alu_a_mux_output_21(\ALUAMUX|alu_a_mux_output[21]~64_combout ),
	.alu_b_mux_output_15(\ALUBMUX|alu_b_mux_output[15]~11_combout ),
	.temp_imemload_output_15(\IDEX|temp_imemload_output [15]),
	.alu_b_mux_output_12(\ALUBMUX|alu_b_mux_output[12]~13_combout ),
	.temp_imemload_output_12(\IDEX|temp_imemload_output [12]),
	.alu_b_mux_output_27(\ALUBMUX|alu_b_mux_output[27]~16_combout ),
	.alu_b_mux_output_18(\ALUBMUX|alu_b_mux_output[18]~18_combout ),
	.alu_b_mux_output_17(\ALUBMUX|alu_b_mux_output[17]~20_combout ),
	.alu_b_mux_output_16(\ALUBMUX|alu_b_mux_output[16]~22_combout ),
	.alu_b_mux_output_31(\ALUBMUX|alu_b_mux_output[31]~24_combout ),
	.alu_b_mux_output_30(\ALUBMUX|alu_b_mux_output[30]~26_combout ),
	.alu_b_mux_output_29(\ALUBMUX|alu_b_mux_output[29]~28_combout ),
	.alu_b_mux_output_28(\ALUBMUX|alu_b_mux_output[28]~30_combout ),
	.alu_b_mux_output_26(\ALUBMUX|alu_b_mux_output[26]~32_combout ),
	.alu_b_mux_output_25(\ALUBMUX|alu_b_mux_output[25]~34_combout ),
	.alu_b_mux_output_24(\ALUBMUX|alu_b_mux_output[24]~36_combout ),
	.alu_b_mux_output_23(\ALUBMUX|alu_b_mux_output[23]~38_combout ),
	.alu_b_mux_output_22(\ALUBMUX|alu_b_mux_output[22]~40_combout ),
	.alu_b_mux_output_21(\ALUBMUX|alu_b_mux_output[21]~42_combout ),
	.alu_b_mux_output_20(\ALUBMUX|alu_b_mux_output[20]~44_combout ),
	.alu_b_mux_output_19(\ALUBMUX|alu_b_mux_output[19]~46_combout ),
	.temp_imemload_output_14(\IDEX|temp_imemload_output [14]),
	.alu_b_mux_output_10(\ALUBMUX|alu_b_mux_output[10]~48_combout ),
	.alu_b_mux_output_14(\ALUBMUX|alu_b_mux_output[14]~50_combout ),
	.alu_b_mux_output_9(\ALUBMUX|alu_b_mux_output[9]~52_combout ),
	.alu_b_mux_output_8(\ALUBMUX|alu_b_mux_output[8]~54_combout ),
	.alu_b_mux_output_7(\ALUBMUX|alu_b_mux_output[7]~56_combout ),
	.alu_b_mux_output_6(\ALUBMUX|alu_b_mux_output[6]~58_combout ),
	.alu_b_mux_output_5(\ALUBMUX|alu_b_mux_output[5]~60_combout ),
	.temp_imemload_output_5(\IDEX|temp_imemload_output [5]),
	.alu_b_mux_output_13(\ALUBMUX|alu_b_mux_output[13]~62_combout ),
	.temp_imemload_output_13(\IDEX|temp_imemload_output [13]),
	.alu_b_mux_output_111(\ALUBMUX|alu_b_mux_output[11]~64_combout ),
	.temp_imemload_output_11(\IDEX|temp_imemload_output [11]),
	.temp_ALUop_output_3(\IDEX|temp_ALUop_output [3]),
	.Mux30(\ALU|Mux30~4_combout ),
	.temp_iMemLoad_31(\EXMEM|temp_iMemLoad [31]),
	.temp_iMemLoad_30(\EXMEM|temp_iMemLoad [30]),
	.temp_iMemLoad_29(\EXMEM|temp_iMemLoad [29]),
	.ex_mem_flush(\HAZARDUNIT|ex_mem_flush~0_combout ),
	.temp_iMemLoad_27(\EXMEM|temp_iMemLoad [27]),
	.temp_iMemLoad_26(\EXMEM|temp_iMemLoad [26]),
	.temp_iMemLoad_28(\EXMEM|temp_iMemLoad [28]),
	.ex_mem_flush1(\HAZARDUNIT|ex_mem_flush~3_combout ),
	.temp_branchSelect1(\EXMEM|temp_branchSelect~q ),
	.ex_mem_flush2(\HAZARDUNIT|ex_mem_flush~4_combout ),
	.ex_mem_flush3(\HAZARDUNIT|ex_mem_flush~5_combout ),
	.wen(\HAZARDUNIT|id_ex_wen~0_combout ),
	.temp_rdat1_1(\EXMEM|temp_rdat1 [1]),
	.temp_npc_1(\EXMEM|temp_npc [1]),
	.temp_pcselect_1(\EXMEM|temp_pcselect [1]),
	.temp_pcselect_0(\EXMEM|temp_pcselect [0]),
	.temp_request_dmemREN_output(\IDEX|temp_request_dmemREN_output~q ),
	.temp_request_dmemWEN_output(\IDEX|temp_request_dmemWEN_output~q ),
	.Mux31(\ALU|Mux31~9_combout ),
	.temp_rdat1_0(\EXMEM|temp_rdat1 [0]),
	.temp_npc_0(\EXMEM|temp_npc [0]),
	.Mux29(\ALU|Mux29~12_combout ),
	.temp_npc_2(\EXMEM|temp_npc [2]),
	.temp_rdat1_2(\EXMEM|temp_rdat1 [2]),
	.Mux28(\ALU|Mux28~6_combout ),
	.temp_npc_3(\EXMEM|temp_npc [3]),
	.temp_rdat1_3(\EXMEM|temp_rdat1 [3]),
	.alu_a_mux_output_32(\ALUAMUX|alu_a_mux_output[3]~65_combout ),
	.Mux26(\ALU|Mux26~6_combout ),
	.temp_npc_5(\EXMEM|temp_npc [5]),
	.temp_npc_4(\EXMEM|temp_npc [4]),
	.temp_rdat1_5(\EXMEM|temp_rdat1 [5]),
	.Mux27(\ALU|Mux27~11_combout ),
	.temp_rdat1_4(\EXMEM|temp_rdat1 [4]),
	.Mux24(\ALU|Mux24~6_combout ),
	.temp_npc_7(\EXMEM|temp_npc [7]),
	.temp_npc_6(\EXMEM|temp_npc [6]),
	.temp_rdat1_7(\EXMEM|temp_rdat1 [7]),
	.Mux25(\ALU|Mux25~6_combout ),
	.temp_rdat1_6(\EXMEM|temp_rdat1 [6]),
	.Mux22(\ALU|Mux22~0_combout ),
	.Mux221(\ALU|Mux22~5_combout ),
	.Mux19(\ALU|Mux19~6_combout ),
	.temp_npc_9(\EXMEM|temp_npc [9]),
	.temp_npc_8(\EXMEM|temp_npc [8]),
	.temp_rdat1_9(\EXMEM|temp_rdat1 [9]),
	.Mux23(\ALU|Mux23~0_combout ),
	.Mux231(\ALU|Mux23~5_combout ),
	.temp_rdat1_8(\EXMEM|temp_rdat1 [8]),
	.Mux20(\ALU|Mux20~0_combout ),
	.Mux201(\ALU|Mux20~5_combout ),
	.temp_npc_11(\EXMEM|temp_npc [11]),
	.temp_npc_10(\EXMEM|temp_npc [10]),
	.temp_rdat1_11(\EXMEM|temp_rdat1 [11]),
	.Mux21(\ALU|Mux21~0_combout ),
	.Mux211(\ALU|Mux21~5_combout ),
	.temp_rdat1_10(\EXMEM|temp_rdat1 [10]),
	.Mux18(\ALU|Mux18~0_combout ),
	.Mux181(\ALU|Mux18~5_combout ),
	.temp_npc_13(\EXMEM|temp_npc [13]),
	.temp_npc_12(\EXMEM|temp_npc [12]),
	.temp_rdat1_13(\EXMEM|temp_rdat1 [13]),
	.Mux191(\ALU|Mux19~7_combout ),
	.Mux192(\ALU|Mux19~12_combout ),
	.temp_rdat1_12(\EXMEM|temp_rdat1 [12]),
	.Mux16(\ALU|Mux16~0_combout ),
	.Mux161(\ALU|Mux16~5_combout ),
	.temp_npc_15(\EXMEM|temp_npc [15]),
	.temp_npc_14(\EXMEM|temp_npc [14]),
	.temp_rdat1_15(\EXMEM|temp_rdat1 [15]),
	.Mux17(\ALU|Mux17~0_combout ),
	.Mux171(\ALU|Mux17~5_combout ),
	.temp_rdat1_14(\EXMEM|temp_rdat1 [14]),
	.Mux14(\ALU|Mux14~0_combout ),
	.Mux141(\ALU|Mux14~4_combout ),
	.temp_npc_17(\EXMEM|temp_npc [17]),
	.temp_npc_16(\EXMEM|temp_npc [16]),
	.temp_rdat1_17(\EXMEM|temp_rdat1 [17]),
	.Mux15(\ALU|Mux15~0_combout ),
	.Mux151(\ALU|Mux15~4_combout ),
	.temp_rdat1_16(\EXMEM|temp_rdat1 [16]),
	.Mux12(\ALU|Mux12~3_combout ),
	.Mux121(\ALU|Mux12~8_combout ),
	.temp_signZero_16(\EXMEM|temp_signZero [16]),
	.temp_npc_19(\EXMEM|temp_npc [19]),
	.temp_npc_18(\EXMEM|temp_npc [18]),
	.temp_rdat1_19(\EXMEM|temp_rdat1 [19]),
	.temp_iMemLoad_17(\EXMEM|temp_iMemLoad [17]),
	.Mux13(\ALU|Mux13~0_combout ),
	.Mux131(\ALU|Mux13~5_combout ),
	.temp_rdat1_18(\EXMEM|temp_rdat1 [18]),
	.temp_iMemLoad_16(\EXMEM|temp_iMemLoad [16]),
	.Mux11(\ALU|Mux11~0_combout ),
	.Mux111(\ALU|Mux11~5_combout ),
	.temp_npc_20(\EXMEM|temp_npc [20]),
	.temp_rdat1_20(\EXMEM|temp_rdat1 [20]),
	.temp_iMemLoad_18(\EXMEM|temp_iMemLoad [18]),
	.Mux10(\ALU|Mux10~0_combout ),
	.Mux101(\ALU|Mux10~5_combout ),
	.temp_npc_21(\EXMEM|temp_npc [21]),
	.temp_rdat1_21(\EXMEM|temp_rdat1 [21]),
	.temp_iMemLoad_19(\EXMEM|temp_iMemLoad [19]),
	.Mux8(\ALU|Mux8~0_combout ),
	.Mux81(\ALU|Mux8~5_combout ),
	.temp_npc_23(\EXMEM|temp_npc [23]),
	.temp_npc_22(\EXMEM|temp_npc [22]),
	.temp_rdat1_23(\EXMEM|temp_rdat1 [23]),
	.temp_iMemLoad_21(\EXMEM|temp_iMemLoad [21]),
	.Mux9(\ALU|Mux9~0_combout ),
	.Mux91(\ALU|Mux9~5_combout ),
	.temp_rdat1_22(\EXMEM|temp_rdat1 [22]),
	.temp_iMemLoad_20(\EXMEM|temp_iMemLoad [20]),
	.Mux6(\ALU|Mux6~7_combout ),
	.temp_npc_25(\EXMEM|temp_npc [25]),
	.temp_npc_24(\EXMEM|temp_npc [24]),
	.temp_rdat1_25(\EXMEM|temp_rdat1 [25]),
	.temp_iMemLoad_23(\EXMEM|temp_iMemLoad [23]),
	.temp_rdat1_24(\EXMEM|temp_rdat1 [24]),
	.temp_iMemLoad_22(\EXMEM|temp_iMemLoad [22]),
	.temp_npc_26(\EXMEM|temp_npc [26]),
	.temp_rdat1_26(\EXMEM|temp_rdat1 [26]),
	.Mux4(\ALU|Mux4~7_combout ),
	.temp_npc_27(\EXMEM|temp_npc [27]),
	.temp_rdat1_27(\EXMEM|temp_rdat1 [27]),
	.Mux2(\ALU|Mux2~14_combout ),
	.temp_npc_29(\EXMEM|temp_npc [29]),
	.temp_npc_28(\EXMEM|temp_npc [28]),
	.temp_rdat1_29(\EXMEM|temp_rdat1 [29]),
	.Mux3(\ALU|Mux3~9_combout ),
	.temp_rdat1_28(\EXMEM|temp_rdat1 [28]),
	.Mux0(\ALU|Mux0~0_combout ),
	.Mux01(\ALU|Mux0~7_combout ),
	.temp_rdat1_31(\EXMEM|temp_rdat1 [31]),
	.temp_npc_31(\EXMEM|temp_npc [31]),
	.temp_npc_30(\EXMEM|temp_npc [30]),
	.Mux1(\ALU|Mux1~2_combout ),
	.temp_rdat1_30(\EXMEM|temp_rdat1 [30]),
	.temp_rdat2_1(temp_rdat2_1),
	.temp_rdat2_2(temp_rdat2_2),
	.temp_rdat2_3(temp_rdat2_3),
	.temp_rdat2_4(temp_rdat2_4),
	.temp_rdat2_5(temp_rdat2_5),
	.temp_rdat2_6(temp_rdat2_6),
	.temp_rdat2_7(temp_rdat2_7),
	.temp_rdat2_8(temp_rdat2_8),
	.temp_rdat2_9(temp_rdat2_9),
	.temp_rdat2_10(temp_rdat2_10),
	.temp_rdat2_11(temp_rdat2_11),
	.temp_rdat2_12(temp_rdat2_12),
	.temp_rdat2_13(temp_rdat2_13),
	.temp_rdat2_14(temp_rdat2_14),
	.temp_rdat2_15(temp_rdat2_15),
	.temp_rdat2_16(temp_rdat2_16),
	.temp_rdat2_17(temp_rdat2_17),
	.temp_rdat2_18(temp_rdat2_18),
	.temp_rdat2_19(temp_rdat2_19),
	.temp_rdat2_20(temp_rdat2_20),
	.temp_rdat2_21(temp_rdat2_21),
	.temp_rdat2_22(temp_rdat2_22),
	.temp_rdat2_23(temp_rdat2_23),
	.temp_rdat2_24(temp_rdat2_24),
	.temp_rdat2_25(temp_rdat2_25),
	.temp_rdat2_26(temp_rdat2_26),
	.temp_rdat2_27(temp_rdat2_27),
	.temp_rdat2_28(temp_rdat2_28),
	.temp_rdat2_29(temp_rdat2_29),
	.temp_rdat2_30(temp_rdat2_30),
	.temp_rdat2_31(temp_rdat2_31),
	.temp_regwrite_output(\IDEX|temp_regwrite_output~q ),
	.temp_regdst_output_1(\IDEX|temp_regdst_output [1]),
	.temp_regdst_output_0(\IDEX|temp_regdst_output [0]),
	.temp_memtoreg_output_0(\IDEX|temp_memtoreg_output [0]),
	.temp_memtoreg_output_1(\IDEX|temp_memtoreg_output [1]),
	.temp_imemload_output_31(\IDEX|temp_imemload_output [31]),
	.temp_imemload_output_30(\IDEX|temp_imemload_output [30]),
	.temp_imemload_output_29(\IDEX|temp_imemload_output [29]),
	.temp_imemload_output_27(\IDEX|temp_imemload_output [27]),
	.temp_imemload_output_26(\IDEX|temp_imemload_output [26]),
	.temp_imemload_output_28(\IDEX|temp_imemload_output [28]),
	.temp_branch_output(\IDEX|temp_branch_output~q ),
	.Equal0(\ALU|Equal0~22_combout ),
	.temp_NPC_output_1(\IDEX|temp_NPC_output [1]),
	.temp_pcselect_output_1(\IDEX|temp_pcselect_output [1]),
	.temp_pcselect_output_0(\IDEX|temp_pcselect_output [0]),
	.temp_NPC_output_0(\IDEX|temp_NPC_output [0]),
	.temp_NPC_output_2(\IDEX|temp_NPC_output [2]),
	.temp_NPC_output_3(\IDEX|temp_NPC_output [3]),
	.temp_NPC_output_5(\IDEX|temp_NPC_output [5]),
	.temp_NPC_output_4(\IDEX|temp_NPC_output [4]),
	.temp_NPC_output_7(\IDEX|temp_NPC_output [7]),
	.temp_NPC_output_6(\IDEX|temp_NPC_output [6]),
	.temp_NPC_output_9(\IDEX|temp_NPC_output [9]),
	.temp_NPC_output_8(\IDEX|temp_NPC_output [8]),
	.temp_NPC_output_11(\IDEX|temp_NPC_output [11]),
	.temp_NPC_output_10(\IDEX|temp_NPC_output [10]),
	.temp_NPC_output_13(\IDEX|temp_NPC_output [13]),
	.temp_NPC_output_12(\IDEX|temp_NPC_output [12]),
	.temp_NPC_output_15(\IDEX|temp_NPC_output [15]),
	.temp_NPC_output_14(\IDEX|temp_NPC_output [14]),
	.temp_NPC_output_17(\IDEX|temp_NPC_output [17]),
	.temp_NPC_output_16(\IDEX|temp_NPC_output [16]),
	.temp_NPC_output_19(\IDEX|temp_NPC_output [19]),
	.temp_NPC_output_18(\IDEX|temp_NPC_output [18]),
	.temp_NPC_output_20(\IDEX|temp_NPC_output [20]),
	.temp_NPC_output_21(\IDEX|temp_NPC_output [21]),
	.temp_NPC_output_23(\IDEX|temp_NPC_output [23]),
	.temp_NPC_output_22(\IDEX|temp_NPC_output [22]),
	.temp_NPC_output_25(\IDEX|temp_NPC_output [25]),
	.temp_NPC_output_24(\IDEX|temp_NPC_output [24]),
	.temp_NPC_output_26(\IDEX|temp_NPC_output [26]),
	.temp_NPC_output_27(\IDEX|temp_NPC_output [27]),
	.temp_NPC_output_29(\IDEX|temp_NPC_output [29]),
	.temp_NPC_output_28(\IDEX|temp_NPC_output [28]),
	.temp_NPC_output_31(\IDEX|temp_NPC_output [31]),
	.temp_NPC_output_30(\IDEX|temp_NPC_output [30]),
	.Mux110(\ALU|Mux1~10_combout ),
	.Mux5(\ALU|Mux5~8_combout ),
	.Mux7(\ALU|Mux7~7_combout ),
	.CLK(CPUCLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

id_ex_latch IDEX(
	.temp_signzerovalue_output_16(\IDEX|temp_signzerovalue_output [16]),
	.temp_halt_out_output1(\IDEX|temp_halt_out_output~q ),
	.temp_ALUop_output_0(\IDEX|temp_ALUop_output [0]),
	.temp_imemload_output_1(\IDEX|temp_imemload_output [1]),
	.temp_imemload_output_7(\IDEX|temp_imemload_output [7]),
	.temp_ALUsrc_output_1(\IDEX|temp_ALUsrc_output [1]),
	.temp_ALUsrc_output_0(\IDEX|temp_ALUsrc_output [0]),
	.temp_rdat_two_output_1(\IDEX|temp_rdat_two_output [1]),
	.temp_imemload_output_17(\IDEX|temp_imemload_output [17]),
	.temp_imemload_output_16(\IDEX|temp_imemload_output [16]),
	.temp_imemload_output_18(\IDEX|temp_imemload_output [18]),
	.temp_imemload_output_19(\IDEX|temp_imemload_output [19]),
	.temp_imemload_output_20(\IDEX|temp_imemload_output [20]),
	.temp_imemload_output_22(\IDEX|temp_imemload_output [22]),
	.temp_imemload_output_21(\IDEX|temp_imemload_output [21]),
	.temp_imemload_output_23(\IDEX|temp_imemload_output [23]),
	.temp_imemload_output_24(\IDEX|temp_imemload_output [24]),
	.temp_imemload_output_25(\IDEX|temp_imemload_output [25]),
	.temp_rdat_one_output_1(\IDEX|temp_rdat_one_output [1]),
	.temp_ALUop_output_1(\IDEX|temp_ALUop_output [1]),
	.temp_imemload_output_0(\IDEX|temp_imemload_output [0]),
	.temp_imemload_output_6(\IDEX|temp_imemload_output [6]),
	.temp_rdat_two_output_0(\IDEX|temp_rdat_two_output [0]),
	.temp_rdat_one_output_0(\IDEX|temp_rdat_one_output [0]),
	.temp_rdat_one_output_2(\IDEX|temp_rdat_one_output [2]),
	.temp_rdat_one_output_4(\IDEX|temp_rdat_one_output [4]),
	.temp_rdat_one_output_3(\IDEX|temp_rdat_one_output [3]),
	.temp_imemload_output_2(\IDEX|temp_imemload_output [2]),
	.temp_imemload_output_8(\IDEX|temp_imemload_output [8]),
	.temp_rdat_two_output_2(\IDEX|temp_rdat_two_output [2]),
	.temp_rdat_one_output_8(\IDEX|temp_rdat_one_output [8]),
	.temp_rdat_one_output_7(\IDEX|temp_rdat_one_output [7]),
	.temp_rdat_one_output_6(\IDEX|temp_rdat_one_output [6]),
	.temp_rdat_one_output_5(\IDEX|temp_rdat_one_output [5]),
	.temp_imemload_output_3(\IDEX|temp_imemload_output [3]),
	.temp_imemload_output_9(\IDEX|temp_imemload_output [9]),
	.temp_rdat_two_output_3(\IDEX|temp_rdat_two_output [3]),
	.temp_rdat_one_output_16(\IDEX|temp_rdat_one_output [16]),
	.temp_rdat_one_output_14(\IDEX|temp_rdat_one_output [14]),
	.temp_rdat_one_output_15(\IDEX|temp_rdat_one_output [15]),
	.temp_rdat_one_output_13(\IDEX|temp_rdat_one_output [13]),
	.temp_rdat_one_output_12(\IDEX|temp_rdat_one_output [12]),
	.temp_rdat_one_output_10(\IDEX|temp_rdat_one_output [10]),
	.temp_rdat_one_output_11(\IDEX|temp_rdat_one_output [11]),
	.temp_rdat_one_output_9(\IDEX|temp_rdat_one_output [9]),
	.temp_imemload_output_4(\IDEX|temp_imemload_output [4]),
	.temp_imemload_output_10(\IDEX|temp_imemload_output [10]),
	.temp_rdat_two_output_4(\IDEX|temp_rdat_two_output [4]),
	.temp_rdat_one_output_31(\IDEX|temp_rdat_one_output [31]),
	.temp_rdat_one_output_30(\IDEX|temp_rdat_one_output [30]),
	.temp_rdat_one_output_29(\IDEX|temp_rdat_one_output [29]),
	.temp_rdat_one_output_26(\IDEX|temp_rdat_one_output [26]),
	.temp_rdat_one_output_25(\IDEX|temp_rdat_one_output [25]),
	.temp_rdat_one_output_28(\IDEX|temp_rdat_one_output [28]),
	.temp_rdat_one_output_27(\IDEX|temp_rdat_one_output [27]),
	.temp_rdat_one_output_17(\IDEX|temp_rdat_one_output [17]),
	.temp_rdat_one_output_20(\IDEX|temp_rdat_one_output [20]),
	.temp_rdat_one_output_19(\IDEX|temp_rdat_one_output [19]),
	.temp_rdat_one_output_18(\IDEX|temp_rdat_one_output [18]),
	.temp_rdat_one_output_24(\IDEX|temp_rdat_one_output [24]),
	.temp_rdat_one_output_23(\IDEX|temp_rdat_one_output [23]),
	.temp_rdat_one_output_22(\IDEX|temp_rdat_one_output [22]),
	.temp_rdat_one_output_21(\IDEX|temp_rdat_one_output [21]),
	.temp_rdat_two_output_15(\IDEX|temp_rdat_two_output [15]),
	.temp_imemload_output_15(\IDEX|temp_imemload_output [15]),
	.temp_rdat_two_output_12(\IDEX|temp_rdat_two_output [12]),
	.temp_imemload_output_12(\IDEX|temp_imemload_output [12]),
	.temp_rdat_two_output_27(\IDEX|temp_rdat_two_output [27]),
	.temp_rdat_two_output_18(\IDEX|temp_rdat_two_output [18]),
	.temp_rdat_two_output_17(\IDEX|temp_rdat_two_output [17]),
	.temp_rdat_two_output_16(\IDEX|temp_rdat_two_output [16]),
	.temp_rdat_two_output_31(\IDEX|temp_rdat_two_output [31]),
	.temp_rdat_two_output_30(\IDEX|temp_rdat_two_output [30]),
	.temp_rdat_two_output_29(\IDEX|temp_rdat_two_output [29]),
	.temp_rdat_two_output_28(\IDEX|temp_rdat_two_output [28]),
	.temp_rdat_two_output_26(\IDEX|temp_rdat_two_output [26]),
	.temp_rdat_two_output_25(\IDEX|temp_rdat_two_output [25]),
	.temp_rdat_two_output_24(\IDEX|temp_rdat_two_output [24]),
	.temp_rdat_two_output_23(\IDEX|temp_rdat_two_output [23]),
	.temp_rdat_two_output_22(\IDEX|temp_rdat_two_output [22]),
	.temp_rdat_two_output_21(\IDEX|temp_rdat_two_output [21]),
	.temp_rdat_two_output_20(\IDEX|temp_rdat_two_output [20]),
	.temp_rdat_two_output_19(\IDEX|temp_rdat_two_output [19]),
	.temp_imemload_output_14(\IDEX|temp_imemload_output [14]),
	.temp_rdat_two_output_10(\IDEX|temp_rdat_two_output [10]),
	.temp_rdat_two_output_14(\IDEX|temp_rdat_two_output [14]),
	.temp_rdat_two_output_9(\IDEX|temp_rdat_two_output [9]),
	.temp_rdat_two_output_8(\IDEX|temp_rdat_two_output [8]),
	.temp_rdat_two_output_7(\IDEX|temp_rdat_two_output [7]),
	.temp_rdat_two_output_6(\IDEX|temp_rdat_two_output [6]),
	.temp_rdat_two_output_5(\IDEX|temp_rdat_two_output [5]),
	.temp_imemload_output_5(\IDEX|temp_imemload_output [5]),
	.temp_rdat_two_output_13(\IDEX|temp_rdat_two_output [13]),
	.temp_imemload_output_13(\IDEX|temp_imemload_output [13]),
	.temp_rdat_two_output_11(\IDEX|temp_rdat_two_output [11]),
	.temp_imemload_output_11(\IDEX|temp_imemload_output [11]),
	.temp_ALUop_output_2(\IDEX|temp_ALUop_output [2]),
	.temp_ALUop_output_3(\IDEX|temp_ALUop_output [3]),
	.ex_mem_flush(\HAZARDUNIT|ex_mem_flush~5_combout ),
	.wen(\HAZARDUNIT|id_ex_wen~0_combout ),
	.temp_request_dmemREN_output1(\IDEX|temp_request_dmemREN_output~q ),
	.temp_imemload_output_171(\IFID|temp_imemload_output [17]),
	.temp_imemload_output_161(\IFID|temp_imemload_output [16]),
	.temp_imemload_output_191(\IFID|temp_imemload_output [19]),
	.temp_imemload_output_181(\IFID|temp_imemload_output [18]),
	.temp_imemload_output_201(\IFID|temp_imemload_output [20]),
	.temp_imemload_output_221(\IFID|temp_imemload_output [22]),
	.temp_imemload_output_211(\IFID|temp_imemload_output [21]),
	.temp_imemload_output_241(\IFID|temp_imemload_output [24]),
	.temp_imemload_output_231(\IFID|temp_imemload_output [23]),
	.temp_imemload_output_251(\IFID|temp_imemload_output [25]),
	.use_after_load(\HAZARDUNIT|use_after_load~6_combout ),
	.temp_request_dmemWEN_output1(\IDEX|temp_request_dmemWEN_output~q ),
	.temp_imemload_output_29(\IFID|temp_imemload_output [29]),
	.temp_imemload_output_31(\IFID|temp_imemload_output [31]),
	.temp_imemload_output_30(\IFID|temp_imemload_output [30]),
	.temp_imemload_output_28(\IFID|temp_imemload_output [28]),
	.Equal3(\CONTROLUNIT|Equal3~0_combout ),
	.temp_imemload_output_27(\IFID|temp_imemload_output [27]),
	.temp_imemload_output_26(\IFID|temp_imemload_output [26]),
	.temp_branch_output1(\IDEX|temp_branch_output~0_combout ),
	.temp_imemload_output_01(\IFID|temp_imemload_output [0]),
	.temp_imemload_output_210(\IFID|temp_imemload_output [2]),
	.temp_imemload_output_32(\IFID|temp_imemload_output [3]),
	.temp_imemload_output_51(\IFID|temp_imemload_output [5]),
	.Equal31(\CONTROLUNIT|Equal3~1_combout ),
	.temp_imemload_output_151(\IFID|temp_imemload_output [15]),
	.temp_imemload_output_141(\IFID|temp_imemload_output [14]),
	.temp_imemload_output_131(\IFID|temp_imemload_output [13]),
	.temp_imemload_output_121(\IFID|temp_imemload_output [12]),
	.temp_imemload_output_111(\IFID|temp_imemload_output [11]),
	.temp_imemload_output_101(\IFID|temp_imemload_output [10]),
	.temp_imemload_output_91(\IFID|temp_imemload_output [9]),
	.temp_imemload_output_81(\IFID|temp_imemload_output [8]),
	.temp_imemload_output_71(\IFID|temp_imemload_output [7]),
	.temp_imemload_output_61(\IFID|temp_imemload_output [6]),
	.temp_imemload_output_110(\IFID|temp_imemload_output [1]),
	.temp_imemload_output_41(\IFID|temp_imemload_output [4]),
	.Equal32(\CONTROLUNIT|Equal3~9_combout ),
	.extended_imm_16(\EXTENDER|extended_imm[16]~0_combout ),
	.WideOr8(\CONTROLUNIT|WideOr8~0_combout ),
	.WideOr2(\CONTROLUNIT|WideOr2~0_combout ),
	.id_ex_flush(\HAZARDUNIT|id_ex_flush~combout ),
	.WideOr4(\CONTROLUNIT|WideOr4~0_combout ),
	.temp_ALUsrc_output(\IDEX|temp_ALUsrc_output~3_combout ),
	.Mux62(\REGISTER|Mux62~9_combout ),
	.Mux621(\REGISTER|Mux62~19_combout ),
	.temp_regwrite_output1(\IDEX|temp_regwrite_output~q ),
	.temp_regdst_output_1(\IDEX|temp_regdst_output [1]),
	.temp_regdst_output_0(\IDEX|temp_regdst_output [0]),
	.temp_memtoreg_output_0(\IDEX|temp_memtoreg_output [0]),
	.temp_memtoreg_output_1(\IDEX|temp_memtoreg_output [1]),
	.Mux30(\REGISTER|Mux30~9_combout ),
	.Mux301(\REGISTER|Mux30~19_combout ),
	.WideOr7(\CONTROLUNIT|WideOr7~0_combout ),
	.WideOr1(\CONTROLUNIT|WideOr1~0_combout ),
	.Mux63(\REGISTER|Mux63~9_combout ),
	.Mux631(\REGISTER|Mux63~19_combout ),
	.Mux31(\REGISTER|Mux31~9_combout ),
	.Mux311(\REGISTER|Mux31~19_combout ),
	.Mux29(\REGISTER|Mux29~9_combout ),
	.Mux291(\REGISTER|Mux29~19_combout ),
	.Mux27(\REGISTER|Mux27~9_combout ),
	.Mux271(\REGISTER|Mux27~19_combout ),
	.Mux28(\REGISTER|Mux28~9_combout ),
	.Mux281(\REGISTER|Mux28~19_combout ),
	.Mux61(\REGISTER|Mux61~9_combout ),
	.Mux611(\REGISTER|Mux61~19_combout ),
	.Mux23(\REGISTER|Mux23~9_combout ),
	.Mux231(\REGISTER|Mux23~19_combout ),
	.Mux24(\REGISTER|Mux24~9_combout ),
	.Mux241(\REGISTER|Mux24~19_combout ),
	.Mux25(\REGISTER|Mux25~9_combout ),
	.Mux251(\REGISTER|Mux25~19_combout ),
	.Mux26(\REGISTER|Mux26~9_combout ),
	.Mux261(\REGISTER|Mux26~19_combout ),
	.Mux60(\REGISTER|Mux60~9_combout ),
	.Mux601(\REGISTER|Mux60~19_combout ),
	.Mux15(\REGISTER|Mux15~9_combout ),
	.Mux151(\REGISTER|Mux15~19_combout ),
	.Mux17(\REGISTER|Mux17~9_combout ),
	.Mux171(\REGISTER|Mux17~19_combout ),
	.Mux16(\REGISTER|Mux16~9_combout ),
	.Mux161(\REGISTER|Mux16~19_combout ),
	.Mux18(\REGISTER|Mux18~9_combout ),
	.Mux181(\REGISTER|Mux18~19_combout ),
	.Mux19(\REGISTER|Mux19~9_combout ),
	.Mux191(\REGISTER|Mux19~19_combout ),
	.Mux21(\REGISTER|Mux21~9_combout ),
	.Mux211(\REGISTER|Mux21~19_combout ),
	.Mux20(\REGISTER|Mux20~9_combout ),
	.Mux201(\REGISTER|Mux20~19_combout ),
	.Mux22(\REGISTER|Mux22~9_combout ),
	.Mux221(\REGISTER|Mux22~19_combout ),
	.Mux59(\REGISTER|Mux59~9_combout ),
	.Mux591(\REGISTER|Mux59~19_combout ),
	.Mux0(\REGISTER|Mux0~9_combout ),
	.Mux01(\REGISTER|Mux0~19_combout ),
	.Mux1(\REGISTER|Mux1~9_combout ),
	.Mux11(\REGISTER|Mux1~19_combout ),
	.Mux2(\REGISTER|Mux2~9_combout ),
	.Mux210(\REGISTER|Mux2~19_combout ),
	.Mux5(\REGISTER|Mux5~9_combout ),
	.Mux51(\REGISTER|Mux5~19_combout ),
	.Mux6(\REGISTER|Mux6~9_combout ),
	.Mux64(\REGISTER|Mux6~19_combout ),
	.Mux3(\REGISTER|Mux3~9_combout ),
	.Mux32(\REGISTER|Mux3~19_combout ),
	.Mux4(\REGISTER|Mux4~9_combout ),
	.Mux41(\REGISTER|Mux4~19_combout ),
	.Mux14(\REGISTER|Mux14~9_combout ),
	.Mux141(\REGISTER|Mux14~19_combout ),
	.Mux111(\REGISTER|Mux11~9_combout ),
	.Mux112(\REGISTER|Mux11~19_combout ),
	.Mux12(\REGISTER|Mux12~9_combout ),
	.Mux121(\REGISTER|Mux12~19_combout ),
	.Mux13(\REGISTER|Mux13~9_combout ),
	.Mux131(\REGISTER|Mux13~19_combout ),
	.Mux7(\REGISTER|Mux7~9_combout ),
	.Mux71(\REGISTER|Mux7~19_combout ),
	.Mux8(\REGISTER|Mux8~9_combout ),
	.Mux81(\REGISTER|Mux8~19_combout ),
	.Mux9(\REGISTER|Mux9~9_combout ),
	.Mux91(\REGISTER|Mux9~19_combout ),
	.Mux10(\REGISTER|Mux10~9_combout ),
	.Mux101(\REGISTER|Mux10~19_combout ),
	.Mux48(\REGISTER|Mux48~9_combout ),
	.Mux481(\REGISTER|Mux48~19_combout ),
	.Mux511(\REGISTER|Mux51~9_combout ),
	.Mux512(\REGISTER|Mux51~19_combout ),
	.Mux36(\REGISTER|Mux36~9_combout ),
	.Mux361(\REGISTER|Mux36~19_combout ),
	.extended_imm_161(\EXTENDER|extended_imm[16]~2_combout ),
	.Mux45(\REGISTER|Mux45~9_combout ),
	.Mux451(\REGISTER|Mux45~19_combout ),
	.Mux46(\REGISTER|Mux46~9_combout ),
	.Mux461(\REGISTER|Mux46~19_combout ),
	.Mux47(\REGISTER|Mux47~9_combout ),
	.Mux471(\REGISTER|Mux47~19_combout ),
	.Mux321(\REGISTER|Mux32~9_combout ),
	.Mux322(\REGISTER|Mux32~19_combout ),
	.Mux33(\REGISTER|Mux33~9_combout ),
	.Mux331(\REGISTER|Mux33~19_combout ),
	.Mux34(\REGISTER|Mux34~9_combout ),
	.Mux341(\REGISTER|Mux34~19_combout ),
	.Mux35(\REGISTER|Mux35~9_combout ),
	.Mux351(\REGISTER|Mux35~19_combout ),
	.Mux37(\REGISTER|Mux37~9_combout ),
	.Mux371(\REGISTER|Mux37~19_combout ),
	.Mux38(\REGISTER|Mux38~9_combout ),
	.Mux381(\REGISTER|Mux38~19_combout ),
	.Mux39(\REGISTER|Mux39~9_combout ),
	.Mux391(\REGISTER|Mux39~19_combout ),
	.Mux40(\REGISTER|Mux40~9_combout ),
	.Mux401(\REGISTER|Mux40~19_combout ),
	.Mux411(\REGISTER|Mux41~9_combout ),
	.Mux412(\REGISTER|Mux41~19_combout ),
	.Mux42(\REGISTER|Mux42~9_combout ),
	.Mux421(\REGISTER|Mux42~19_combout ),
	.Mux43(\REGISTER|Mux43~9_combout ),
	.Mux431(\REGISTER|Mux43~19_combout ),
	.Mux44(\REGISTER|Mux44~9_combout ),
	.Mux441(\REGISTER|Mux44~19_combout ),
	.Mux53(\REGISTER|Mux53~9_combout ),
	.Mux531(\REGISTER|Mux53~19_combout ),
	.Mux49(\REGISTER|Mux49~9_combout ),
	.Mux491(\REGISTER|Mux49~19_combout ),
	.Mux54(\REGISTER|Mux54~9_combout ),
	.Mux541(\REGISTER|Mux54~19_combout ),
	.Mux55(\REGISTER|Mux55~9_combout ),
	.Mux551(\REGISTER|Mux55~19_combout ),
	.Mux56(\REGISTER|Mux56~9_combout ),
	.Mux561(\REGISTER|Mux56~19_combout ),
	.Mux57(\REGISTER|Mux57~9_combout ),
	.Mux571(\REGISTER|Mux57~19_combout ),
	.Mux58(\REGISTER|Mux58~9_combout ),
	.Mux581(\REGISTER|Mux58~19_combout ),
	.Mux50(\REGISTER|Mux50~9_combout ),
	.Mux501(\REGISTER|Mux50~19_combout ),
	.Mux52(\REGISTER|Mux52~9_combout ),
	.Mux521(\REGISTER|Mux52~19_combout ),
	.WideOr6(\CONTROLUNIT|WideOr6~0_combout ),
	.WideOr0(\CONTROLUNIT|WideOr0~0_combout ),
	.halt_out(\CONTROLUNIT|halt_out~0_combout ),
	.temp_imemload_output_311(\IDEX|temp_imemload_output [31]),
	.temp_imemload_output_301(\IDEX|temp_imemload_output [30]),
	.temp_imemload_output_291(\IDEX|temp_imemload_output [29]),
	.temp_imemload_output_271(\IDEX|temp_imemload_output [27]),
	.temp_imemload_output_261(\IDEX|temp_imemload_output [26]),
	.temp_imemload_output_281(\IDEX|temp_imemload_output [28]),
	.temp_branch_output2(\IDEX|temp_branch_output~q ),
	.temp_NPC_output_1(\IDEX|temp_NPC_output [1]),
	.temp_pcselect_output_1(\IDEX|temp_pcselect_output [1]),
	.temp_pcselect_output_0(\IDEX|temp_pcselect_output [0]),
	.temp_NPC_output_0(\IDEX|temp_NPC_output [0]),
	.temp_NPC_output_2(\IDEX|temp_NPC_output [2]),
	.temp_NPC_output_3(\IDEX|temp_NPC_output [3]),
	.temp_NPC_output_5(\IDEX|temp_NPC_output [5]),
	.temp_NPC_output_4(\IDEX|temp_NPC_output [4]),
	.temp_NPC_output_7(\IDEX|temp_NPC_output [7]),
	.temp_NPC_output_6(\IDEX|temp_NPC_output [6]),
	.temp_NPC_output_9(\IDEX|temp_NPC_output [9]),
	.temp_NPC_output_8(\IDEX|temp_NPC_output [8]),
	.temp_NPC_output_11(\IDEX|temp_NPC_output [11]),
	.temp_NPC_output_10(\IDEX|temp_NPC_output [10]),
	.temp_NPC_output_13(\IDEX|temp_NPC_output [13]),
	.temp_NPC_output_12(\IDEX|temp_NPC_output [12]),
	.temp_NPC_output_15(\IDEX|temp_NPC_output [15]),
	.temp_NPC_output_14(\IDEX|temp_NPC_output [14]),
	.temp_NPC_output_17(\IDEX|temp_NPC_output [17]),
	.temp_NPC_output_16(\IDEX|temp_NPC_output [16]),
	.temp_NPC_output_19(\IDEX|temp_NPC_output [19]),
	.temp_NPC_output_18(\IDEX|temp_NPC_output [18]),
	.temp_NPC_output_20(\IDEX|temp_NPC_output [20]),
	.temp_NPC_output_21(\IDEX|temp_NPC_output [21]),
	.temp_NPC_output_23(\IDEX|temp_NPC_output [23]),
	.temp_NPC_output_22(\IDEX|temp_NPC_output [22]),
	.temp_NPC_output_25(\IDEX|temp_NPC_output [25]),
	.temp_NPC_output_24(\IDEX|temp_NPC_output [24]),
	.temp_NPC_output_26(\IDEX|temp_NPC_output [26]),
	.temp_NPC_output_27(\IDEX|temp_NPC_output [27]),
	.temp_NPC_output_29(\IDEX|temp_NPC_output [29]),
	.temp_NPC_output_28(\IDEX|temp_NPC_output [28]),
	.temp_NPC_output_31(\IDEX|temp_NPC_output [31]),
	.temp_NPC_output_30(\IDEX|temp_NPC_output [30]),
	.halt_out1(\CONTROLUNIT|halt_out~3_combout ),
	.WideOr3(\CONTROLUNIT|WideOr3~0_combout ),
	.WideOr10(\CONTROLUNIT|WideOr10~0_combout ),
	.memtoreg(\CONTROLUNIT|memtoreg~0_combout ),
	.temp_NPC_output_110(\IFID|temp_NPC_output [1]),
	.WideOr9(\CONTROLUNIT|WideOr9~0_combout ),
	.temp_NPC_output_01(\IFID|temp_NPC_output [0]),
	.temp_NPC_output_210(\IFID|temp_NPC_output [2]),
	.temp_NPC_output_32(\IFID|temp_NPC_output [3]),
	.temp_NPC_output_51(\IFID|temp_NPC_output [5]),
	.temp_NPC_output_41(\IFID|temp_NPC_output [4]),
	.temp_NPC_output_71(\IFID|temp_NPC_output [7]),
	.temp_NPC_output_61(\IFID|temp_NPC_output [6]),
	.temp_NPC_output_91(\IFID|temp_NPC_output [9]),
	.temp_NPC_output_81(\IFID|temp_NPC_output [8]),
	.temp_NPC_output_111(\IFID|temp_NPC_output [11]),
	.temp_NPC_output_101(\IFID|temp_NPC_output [10]),
	.temp_NPC_output_131(\IFID|temp_NPC_output [13]),
	.temp_NPC_output_121(\IFID|temp_NPC_output [12]),
	.temp_NPC_output_151(\IFID|temp_NPC_output [15]),
	.temp_NPC_output_141(\IFID|temp_NPC_output [14]),
	.temp_NPC_output_171(\IFID|temp_NPC_output [17]),
	.temp_NPC_output_161(\IFID|temp_NPC_output [16]),
	.temp_NPC_output_191(\IFID|temp_NPC_output [19]),
	.temp_NPC_output_181(\IFID|temp_NPC_output [18]),
	.temp_NPC_output_201(\IFID|temp_NPC_output [20]),
	.temp_NPC_output_211(\IFID|temp_NPC_output [21]),
	.temp_NPC_output_231(\IFID|temp_NPC_output [23]),
	.temp_NPC_output_221(\IFID|temp_NPC_output [22]),
	.temp_NPC_output_251(\IFID|temp_NPC_output [25]),
	.temp_NPC_output_241(\IFID|temp_NPC_output [24]),
	.temp_NPC_output_261(\IFID|temp_NPC_output [26]),
	.temp_NPC_output_271(\IFID|temp_NPC_output [27]),
	.temp_NPC_output_291(\IFID|temp_NPC_output [29]),
	.temp_NPC_output_281(\IFID|temp_NPC_output [28]),
	.temp_NPC_output_311(\IFID|temp_NPC_output [31]),
	.temp_NPC_output_301(\IFID|temp_NPC_output [30]),
	.CLK(CPUCLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

if_id_latch IFID(
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.ex_mem_flush(\HAZARDUNIT|ex_mem_flush~5_combout ),
	.Mux30(\NPCMUX|Mux30~1_combout ),
	.ccifiwait_0(ccifiwait_0),
	.temp_imemload_output_17(\IFID|temp_imemload_output [17]),
	.temp_imemload_output_16(\IFID|temp_imemload_output [16]),
	.temp_imemload_output_19(\IFID|temp_imemload_output [19]),
	.temp_imemload_output_18(\IFID|temp_imemload_output [18]),
	.temp_imemload_output_20(\IFID|temp_imemload_output [20]),
	.temp_imemload_output_22(\IFID|temp_imemload_output [22]),
	.temp_imemload_output_21(\IFID|temp_imemload_output [21]),
	.temp_imemload_output_24(\IFID|temp_imemload_output [24]),
	.temp_imemload_output_23(\IFID|temp_imemload_output [23]),
	.temp_imemload_output_25(\IFID|temp_imemload_output [25]),
	.Mux31(\NPCMUX|Mux31~2_combout ),
	.Mux29(\NPCMUX|Mux29~1_combout ),
	.Mux28(\NPCMUX|Mux28~1_combout ),
	.Mux26(\NPCMUX|Mux26~1_combout ),
	.Mux27(\NPCMUX|Mux27~1_combout ),
	.Mux24(\NPCMUX|Mux24~1_combout ),
	.Mux25(\NPCMUX|Mux25~1_combout ),
	.Mux22(\NPCMUX|Mux22~1_combout ),
	.Mux23(\NPCMUX|Mux23~1_combout ),
	.Mux20(\NPCMUX|Mux20~1_combout ),
	.Mux21(\NPCMUX|Mux21~1_combout ),
	.Mux18(\NPCMUX|Mux18~1_combout ),
	.Mux19(\NPCMUX|Mux19~1_combout ),
	.Mux16(\NPCMUX|Mux16~1_combout ),
	.Mux17(\NPCMUX|Mux17~1_combout ),
	.Mux14(\NPCMUX|Mux14~1_combout ),
	.Mux15(\NPCMUX|Mux15~1_combout ),
	.Mux12(\NPCMUX|Mux12~1_combout ),
	.Mux13(\NPCMUX|Mux13~1_combout ),
	.Mux11(\NPCMUX|Mux11~1_combout ),
	.Mux10(\NPCMUX|Mux10~1_combout ),
	.Mux8(\NPCMUX|Mux8~1_combout ),
	.Mux9(\NPCMUX|Mux9~1_combout ),
	.Mux6(\NPCMUX|Mux6~1_combout ),
	.Mux7(\NPCMUX|Mux7~1_combout ),
	.Mux5(\NPCMUX|Mux5~1_combout ),
	.Mux4(\NPCMUX|Mux4~1_combout ),
	.Mux2(\NPCMUX|Mux2~1_combout ),
	.Mux3(\NPCMUX|Mux3~3_combout ),
	.Mux0(\NPCMUX|Mux0~1_combout ),
	.Mux1(\NPCMUX|Mux1~1_combout ),
	.temp_imemload_output_29(\IFID|temp_imemload_output [29]),
	.temp_imemload_output_31(\IFID|temp_imemload_output [31]),
	.temp_imemload_output_30(\IFID|temp_imemload_output [30]),
	.temp_imemload_output_28(\IFID|temp_imemload_output [28]),
	.temp_imemload_output_27(\IFID|temp_imemload_output [27]),
	.temp_imemload_output_26(\IFID|temp_imemload_output [26]),
	.temp_imemload_output_0(\IFID|temp_imemload_output [0]),
	.temp_imemload_output_2(\IFID|temp_imemload_output [2]),
	.temp_imemload_output_3(\IFID|temp_imemload_output [3]),
	.temp_imemload_output_5(\IFID|temp_imemload_output [5]),
	.temp_imemload_output_15(\IFID|temp_imemload_output [15]),
	.temp_imemload_output_14(\IFID|temp_imemload_output [14]),
	.temp_imemload_output_13(\IFID|temp_imemload_output [13]),
	.temp_imemload_output_12(\IFID|temp_imemload_output [12]),
	.temp_imemload_output_11(\IFID|temp_imemload_output [11]),
	.temp_imemload_output_10(\IFID|temp_imemload_output [10]),
	.temp_imemload_output_9(\IFID|temp_imemload_output [9]),
	.temp_imemload_output_8(\IFID|temp_imemload_output [8]),
	.temp_imemload_output_7(\IFID|temp_imemload_output [7]),
	.temp_imemload_output_6(\IFID|temp_imemload_output [6]),
	.temp_imemload_output_1(\IFID|temp_imemload_output [1]),
	.temp_imemload_output_4(\IFID|temp_imemload_output [4]),
	.wen(\HAZARDUNIT|pc_wen~3_combout ),
	.temp_NPC_output_1(\IFID|temp_NPC_output [1]),
	.temp_NPC_output_0(\IFID|temp_NPC_output [0]),
	.temp_NPC_output_2(\IFID|temp_NPC_output [2]),
	.temp_NPC_output_3(\IFID|temp_NPC_output [3]),
	.temp_NPC_output_5(\IFID|temp_NPC_output [5]),
	.temp_NPC_output_4(\IFID|temp_NPC_output [4]),
	.temp_NPC_output_7(\IFID|temp_NPC_output [7]),
	.temp_NPC_output_6(\IFID|temp_NPC_output [6]),
	.temp_NPC_output_9(\IFID|temp_NPC_output [9]),
	.temp_NPC_output_8(\IFID|temp_NPC_output [8]),
	.temp_NPC_output_11(\IFID|temp_NPC_output [11]),
	.temp_NPC_output_10(\IFID|temp_NPC_output [10]),
	.temp_NPC_output_13(\IFID|temp_NPC_output [13]),
	.temp_NPC_output_12(\IFID|temp_NPC_output [12]),
	.temp_NPC_output_15(\IFID|temp_NPC_output [15]),
	.temp_NPC_output_14(\IFID|temp_NPC_output [14]),
	.temp_NPC_output_17(\IFID|temp_NPC_output [17]),
	.temp_NPC_output_16(\IFID|temp_NPC_output [16]),
	.temp_NPC_output_19(\IFID|temp_NPC_output [19]),
	.temp_NPC_output_18(\IFID|temp_NPC_output [18]),
	.temp_NPC_output_20(\IFID|temp_NPC_output [20]),
	.temp_NPC_output_21(\IFID|temp_NPC_output [21]),
	.temp_NPC_output_23(\IFID|temp_NPC_output [23]),
	.temp_NPC_output_22(\IFID|temp_NPC_output [22]),
	.temp_NPC_output_25(\IFID|temp_NPC_output [25]),
	.temp_NPC_output_24(\IFID|temp_NPC_output [24]),
	.temp_NPC_output_26(\IFID|temp_NPC_output [26]),
	.temp_NPC_output_27(\IFID|temp_NPC_output [27]),
	.temp_NPC_output_29(\IFID|temp_NPC_output [29]),
	.temp_NPC_output_28(\IFID|temp_NPC_output [28]),
	.temp_NPC_output_31(\IFID|temp_NPC_output [31]),
	.temp_NPC_output_30(\IFID|temp_NPC_output [30]),
	.CLK(CPUCLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

forward FORWADUNIT(
	.temp_branchDest_0(\EXMEM|temp_branchDest [0]),
	.temp_branchDest_4(\EXMEM|temp_branchDest [4]),
	.temp_branchDest_3(\EXMEM|temp_branchDest [3]),
	.temp_branchDest_2(\EXMEM|temp_branchDest [2]),
	.temp_branchDest_1(\EXMEM|temp_branchDest [1]),
	.temp_regwrite(\EXMEM|temp_regwrite~q ),
	.temp_imemload_output_17(\IDEX|temp_imemload_output [17]),
	.temp_imemload_output_16(\IDEX|temp_imemload_output [16]),
	.temp_imemload_output_18(\IDEX|temp_imemload_output [18]),
	.temp_imemload_output_19(\IDEX|temp_imemload_output [19]),
	.temp_imemload_output_20(\IDEX|temp_imemload_output [20]),
	.temp_memtoreg_0(\EXMEM|temp_memtoreg [0]),
	.temp_memtoreg_1(\EXMEM|temp_memtoreg [1]),
	.always0(\FORWADUNIT|always0~7_combout ),
	.temp_regwrite1(\MEMWB|temp_regwrite~q ),
	.always01(\FORWADUNIT|always0~8_combout ),
	.temp_branchDest_11(\MEMWB|temp_branchDest [1]),
	.temp_branchDest_01(\MEMWB|temp_branchDest [0]),
	.temp_branchDest_31(\MEMWB|temp_branchDest [3]),
	.temp_branchDest_21(\MEMWB|temp_branchDest [2]),
	.temp_branchDest_41(\MEMWB|temp_branchDest [4]),
	.always02(\FORWADUNIT|always0~12_combout ),
	.always03(\FORWADUNIT|always0~13_combout ),
	.forwardb_1(\FORWADUNIT|forwardb[1]~0_combout ),
	.temp_imemload_output_22(\IDEX|temp_imemload_output [22]),
	.temp_imemload_output_21(\IDEX|temp_imemload_output [21]),
	.temp_imemload_output_23(\IDEX|temp_imemload_output [23]),
	.temp_imemload_output_24(\IDEX|temp_imemload_output [24]),
	.temp_imemload_output_25(\IDEX|temp_imemload_output [25]),
	.forwarda_1(\FORWADUNIT|forwarda[1]~3_combout ),
	.always04(\FORWADUNIT|always0~16_combout ),
	.always05(\FORWADUNIT|always0~17_combout ),
	.always06(\FORWADUNIT|always0~18_combout ),
	.always07(\FORWADUNIT|always0~19_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

hazard_unit HAZARDUNIT(
	.temp_zeroFlag(\EXMEM|temp_zeroFlag~q ),
	.temp_dmemWEN(temp_dmemWEN),
	.temp_dmemREN(temp_dmemREN),
	.always1(always1),
	.temp_halt_out(\EXMEM|temp_halt_out~q ),
	.temp_imemload_output_17(\IDEX|temp_imemload_output [17]),
	.temp_imemload_output_16(\IDEX|temp_imemload_output [16]),
	.temp_imemload_output_18(\IDEX|temp_imemload_output [18]),
	.temp_imemload_output_19(\IDEX|temp_imemload_output [19]),
	.temp_imemload_output_20(\IDEX|temp_imemload_output [20]),
	.temp_iMemLoad_0(\EXMEM|temp_iMemLoad [0]),
	.temp_iMemLoad_1(\EXMEM|temp_iMemLoad [1]),
	.temp_iMemLoad_4(\EXMEM|temp_iMemLoad [4]),
	.temp_iMemLoad_3(\EXMEM|temp_iMemLoad [3]),
	.temp_iMemLoad_2(\EXMEM|temp_iMemLoad [2]),
	.temp_iMemLoad_5(\EXMEM|temp_iMemLoad [5]),
	.temp_iMemLoad_31(\EXMEM|temp_iMemLoad [31]),
	.temp_iMemLoad_30(\EXMEM|temp_iMemLoad [30]),
	.temp_iMemLoad_29(\EXMEM|temp_iMemLoad [29]),
	.ex_mem_flush(\HAZARDUNIT|ex_mem_flush~0_combout ),
	.temp_iMemLoad_27(\EXMEM|temp_iMemLoad [27]),
	.temp_iMemLoad_26(\EXMEM|temp_iMemLoad [26]),
	.temp_iMemLoad_28(\EXMEM|temp_iMemLoad [28]),
	.ex_mem_flush1(\HAZARDUNIT|ex_mem_flush~3_combout ),
	.temp_branchSelect(\EXMEM|temp_branchSelect~q ),
	.ex_mem_flush2(\HAZARDUNIT|ex_mem_flush~4_combout ),
	.ex_mem_flush3(\HAZARDUNIT|ex_mem_flush~5_combout ),
	.id_ex_wen(\HAZARDUNIT|id_ex_wen~0_combout ),
	.ccifiwait_0(ccifiwait_0),
	.temp_request_dmemREN_output(\IDEX|temp_request_dmemREN_output~q ),
	.temp_imemload_output_171(\IFID|temp_imemload_output [17]),
	.temp_imemload_output_161(\IFID|temp_imemload_output [16]),
	.temp_imemload_output_191(\IFID|temp_imemload_output [19]),
	.temp_imemload_output_181(\IFID|temp_imemload_output [18]),
	.temp_imemload_output_201(\IFID|temp_imemload_output [20]),
	.temp_imemload_output_22(\IFID|temp_imemload_output [22]),
	.temp_imemload_output_21(\IFID|temp_imemload_output [21]),
	.temp_imemload_output_24(\IFID|temp_imemload_output [24]),
	.temp_imemload_output_23(\IFID|temp_imemload_output [23]),
	.temp_imemload_output_25(\IFID|temp_imemload_output [25]),
	.use_after_load(\HAZARDUNIT|use_after_load~6_combout ),
	.pc_wen(\HAZARDUNIT|pc_wen~2_combout ),
	.id_ex_flush1(\HAZARDUNIT|id_ex_flush~combout ),
	.pc_wen1(\HAZARDUNIT|pc_wen~3_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

alu ALU(
	.temp_ALUop_output_0(\IDEX|temp_ALUop_output [0]),
	.temp_imemload_output_7(\IDEX|temp_imemload_output [7]),
	.temp_ALUsrc_output_1(\IDEX|temp_ALUsrc_output [1]),
	.temp_ALUsrc_output_0(\IDEX|temp_ALUsrc_output [0]),
	.Mux30(\alusourceMUX|Mux30~0_combout ),
	.alu_b_mux_output_1(\ALUBMUX|alu_b_mux_output[1]~0_combout ),
	.alu_b_mux_output_11(\ALUBMUX|alu_b_mux_output[1]~1_combout ),
	.Mux16(\alusourceMUX|Mux16~0_combout ),
	.Mux301(\alusourceMUX|Mux30~1_combout ),
	.alu_a_mux_output_1(\ALUAMUX|alu_a_mux_output[1]~1_combout ),
	.temp_ALUop_output_1(\IDEX|temp_ALUop_output [1]),
	.alu_b_mux_output_0(\ALUBMUX|alu_b_mux_output[0]~2_combout ),
	.temp_imemload_output_6(\IDEX|temp_imemload_output [6]),
	.Mux31(\alusourceMUX|Mux31~0_combout ),
	.alu_b_mux_output_01(\ALUBMUX|alu_b_mux_output[0]~3_combout ),
	.alu_a_mux_output_0(\ALUAMUX|alu_a_mux_output[0]~3_combout ),
	.alu_a_mux_output_2(\ALUAMUX|alu_a_mux_output[2]~5_combout ),
	.Mux311(\alusourceMUX|Mux31~1_combout ),
	.alu_a_mux_output_4(\ALUAMUX|alu_a_mux_output[4]~7_combout ),
	.alu_a_mux_output_3(\ALUAMUX|alu_a_mux_output[3]~8_combout ),
	.alu_a_mux_output_31(\ALUAMUX|alu_a_mux_output[3]~9_combout ),
	.Mux29(\alusourceMUX|Mux29~0_combout ),
	.alu_b_mux_output_2(\ALUBMUX|alu_b_mux_output[2]~5_combout ),
	.Mux291(\alusourceMUX|Mux29~1_combout ),
	.alu_a_mux_output_8(\ALUAMUX|alu_a_mux_output[8]~11_combout ),
	.alu_a_mux_output_7(\ALUAMUX|alu_a_mux_output[7]~13_combout ),
	.alu_a_mux_output_6(\ALUAMUX|alu_a_mux_output[6]~15_combout ),
	.alu_a_mux_output_5(\ALUAMUX|alu_a_mux_output[5]~17_combout ),
	.Mux28(\alusourceMUX|Mux28~0_combout ),
	.alu_b_mux_output_3(\ALUBMUX|alu_b_mux_output[3]~7_combout ),
	.Mux281(\alusourceMUX|Mux28~1_combout ),
	.alu_a_mux_output_16(\ALUAMUX|alu_a_mux_output[16]~20_combout ),
	.alu_a_mux_output_14(\ALUAMUX|alu_a_mux_output[14]~22_combout ),
	.alu_a_mux_output_15(\ALUAMUX|alu_a_mux_output[15]~24_combout ),
	.alu_a_mux_output_13(\ALUAMUX|alu_a_mux_output[13]~26_combout ),
	.alu_a_mux_output_12(\ALUAMUX|alu_a_mux_output[12]~28_combout ),
	.alu_a_mux_output_10(\ALUAMUX|alu_a_mux_output[10]~30_combout ),
	.alu_a_mux_output_11(\ALUAMUX|alu_a_mux_output[11]~32_combout ),
	.alu_a_mux_output_9(\ALUAMUX|alu_a_mux_output[9]~34_combout ),
	.Mux27(\alusourceMUX|Mux27~0_combout ),
	.alu_b_mux_output_4(\ALUBMUX|alu_b_mux_output[4]~9_combout ),
	.Mux271(\alusourceMUX|Mux27~1_combout ),
	.alu_a_mux_output_311(\ALUAMUX|alu_a_mux_output[31]~36_combout ),
	.alu_a_mux_output_30(\ALUAMUX|alu_a_mux_output[30]~38_combout ),
	.alu_a_mux_output_29(\ALUAMUX|alu_a_mux_output[29]~40_combout ),
	.alu_a_mux_output_26(\ALUAMUX|alu_a_mux_output[26]~42_combout ),
	.alu_a_mux_output_25(\ALUAMUX|alu_a_mux_output[25]~44_combout ),
	.alu_a_mux_output_28(\ALUAMUX|alu_a_mux_output[28]~46_combout ),
	.alu_a_mux_output_27(\ALUAMUX|alu_a_mux_output[27]~48_combout ),
	.alu_a_mux_output_17(\ALUAMUX|alu_a_mux_output[17]~50_combout ),
	.alu_a_mux_output_20(\ALUAMUX|alu_a_mux_output[20]~52_combout ),
	.alu_a_mux_output_19(\ALUAMUX|alu_a_mux_output[19]~54_combout ),
	.alu_a_mux_output_18(\ALUAMUX|alu_a_mux_output[18]~56_combout ),
	.alu_a_mux_output_24(\ALUAMUX|alu_a_mux_output[24]~58_combout ),
	.alu_a_mux_output_23(\ALUAMUX|alu_a_mux_output[23]~60_combout ),
	.alu_a_mux_output_22(\ALUAMUX|alu_a_mux_output[22]~62_combout ),
	.alu_a_mux_output_21(\ALUAMUX|alu_a_mux_output[21]~64_combout ),
	.Mux161(\alusourceMUX|Mux16~1_combout ),
	.Mux19(\alusourceMUX|Mux19~0_combout ),
	.Mux4(\alusourceMUX|Mux4~0_combout ),
	.Mux13(\alusourceMUX|Mux13~0_combout ),
	.Mux14(\alusourceMUX|Mux14~0_combout ),
	.Mux15(\alusourceMUX|Mux15~0_combout ),
	.Mux0(\alusourceMUX|Mux0~0_combout ),
	.Mux1(\alusourceMUX|Mux1~0_combout ),
	.Mux2(\alusourceMUX|Mux2~0_combout ),
	.Mux3(\alusourceMUX|Mux3~0_combout ),
	.Mux5(\alusourceMUX|Mux5~0_combout ),
	.Mux6(\alusourceMUX|Mux6~0_combout ),
	.Mux7(\alusourceMUX|Mux7~0_combout ),
	.Mux8(\alusourceMUX|Mux8~0_combout ),
	.Mux9(\alusourceMUX|Mux9~0_combout ),
	.Mux10(\alusourceMUX|Mux10~0_combout ),
	.Mux11(\alusourceMUX|Mux11~0_combout ),
	.Mux12(\alusourceMUX|Mux12~0_combout ),
	.Mux17(\alusourceMUX|Mux17~0_combout ),
	.Mux21(\alusourceMUX|Mux21~0_combout ),
	.alu_b_mux_output_14(\ALUBMUX|alu_b_mux_output[14]~50_combout ),
	.Mux22(\alusourceMUX|Mux22~0_combout ),
	.Mux23(\alusourceMUX|Mux23~0_combout ),
	.alu_b_mux_output_7(\ALUBMUX|alu_b_mux_output[7]~56_combout ),
	.Mux24(\alusourceMUX|Mux24~0_combout ),
	.alu_b_mux_output_6(\ALUBMUX|alu_b_mux_output[6]~58_combout ),
	.Mux25(\alusourceMUX|Mux25~0_combout ),
	.alu_b_mux_output_5(\ALUBMUX|alu_b_mux_output[5]~60_combout ),
	.temp_imemload_output_5(\IDEX|temp_imemload_output [5]),
	.Mux26(\alusourceMUX|Mux26~0_combout ),
	.Mux18(\alusourceMUX|Mux18~0_combout ),
	.Mux20(\alusourceMUX|Mux20~0_combout ),
	.temp_ALUop_output_2(\IDEX|temp_ALUop_output [2]),
	.temp_ALUop_output_3(\IDEX|temp_ALUop_output [3]),
	.Mux302(\ALU|Mux30~4_combout ),
	.Mux171(\alusourceMUX|Mux17~1_combout ),
	.Mux312(\ALU|Mux31~9_combout ),
	.Mux292(\ALU|Mux29~12_combout ),
	.Mux282(\ALU|Mux28~6_combout ),
	.alu_a_mux_output_32(\ALUAMUX|alu_a_mux_output[3]~65_combout ),
	.Mux261(\ALU|Mux26~6_combout ),
	.Mux272(\ALU|Mux27~11_combout ),
	.Mux241(\ALU|Mux24~6_combout ),
	.Mux251(\ALU|Mux25~6_combout ),
	.Mux221(\ALU|Mux22~0_combout ),
	.Mux222(\ALU|Mux22~5_combout ),
	.Mux191(\ALU|Mux19~6_combout ),
	.Mux231(\ALU|Mux23~0_combout ),
	.Mux232(\ALU|Mux23~5_combout ),
	.Mux201(\ALU|Mux20~0_combout ),
	.Mux202(\ALU|Mux20~5_combout ),
	.Mux211(\ALU|Mux21~0_combout ),
	.Mux212(\ALU|Mux21~5_combout ),
	.Mux181(\ALU|Mux18~0_combout ),
	.Mux182(\ALU|Mux18~5_combout ),
	.Mux192(\ALU|Mux19~7_combout ),
	.Mux193(\ALU|Mux19~12_combout ),
	.Mux162(\ALU|Mux16~0_combout ),
	.Mux163(\ALU|Mux16~5_combout ),
	.Mux172(\ALU|Mux17~0_combout ),
	.Mux173(\ALU|Mux17~5_combout ),
	.Mux141(\ALU|Mux14~0_combout ),
	.Mux142(\ALU|Mux14~4_combout ),
	.Mux151(\ALU|Mux15~0_combout ),
	.Mux152(\ALU|Mux15~4_combout ),
	.Mux121(\ALU|Mux12~3_combout ),
	.Mux122(\ALU|Mux12~8_combout ),
	.Mux131(\ALU|Mux13~0_combout ),
	.Mux132(\ALU|Mux13~5_combout ),
	.Mux111(\ALU|Mux11~0_combout ),
	.Mux112(\ALU|Mux11~5_combout ),
	.Mux101(\ALU|Mux10~0_combout ),
	.Mux102(\ALU|Mux10~5_combout ),
	.Mux81(\ALU|Mux8~0_combout ),
	.Mux82(\ALU|Mux8~5_combout ),
	.Mux91(\ALU|Mux9~0_combout ),
	.Mux92(\ALU|Mux9~5_combout ),
	.Mux61(\ALU|Mux6~7_combout ),
	.Mux41(\ALU|Mux4~7_combout ),
	.Mux210(\ALU|Mux2~14_combout ),
	.Mux32(\ALU|Mux3~9_combout ),
	.Mux01(\ALU|Mux0~0_combout ),
	.Mux02(\ALU|Mux0~7_combout ),
	.Mux110(\ALU|Mux1~2_combout ),
	.Equal0(\ALU|Equal0~22_combout ),
	.Mux113(\ALU|Mux1~10_combout ),
	.Mux51(\ALU|Mux5~8_combout ),
	.Mux71(\ALU|Mux7~7_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

control_unit CONTROLUNIT(
	.temp_imemload_output_17(\IFID|temp_imemload_output [17]),
	.temp_imemload_output_16(\IFID|temp_imemload_output [16]),
	.temp_imemload_output_19(\IFID|temp_imemload_output [19]),
	.temp_imemload_output_18(\IFID|temp_imemload_output [18]),
	.temp_imemload_output_20(\IFID|temp_imemload_output [20]),
	.temp_imemload_output_22(\IFID|temp_imemload_output [22]),
	.temp_imemload_output_21(\IFID|temp_imemload_output [21]),
	.temp_imemload_output_24(\IFID|temp_imemload_output [24]),
	.temp_imemload_output_23(\IFID|temp_imemload_output [23]),
	.temp_imemload_output_25(\IFID|temp_imemload_output [25]),
	.temp_imemload_output_29(\IFID|temp_imemload_output [29]),
	.temp_imemload_output_31(\IFID|temp_imemload_output [31]),
	.temp_imemload_output_30(\IFID|temp_imemload_output [30]),
	.temp_imemload_output_28(\IFID|temp_imemload_output [28]),
	.Equal3(\CONTROLUNIT|Equal3~0_combout ),
	.temp_imemload_output_27(\IFID|temp_imemload_output [27]),
	.temp_imemload_output_26(\IFID|temp_imemload_output [26]),
	.temp_branch_output(\IDEX|temp_branch_output~0_combout ),
	.temp_imemload_output_0(\IFID|temp_imemload_output [0]),
	.temp_imemload_output_2(\IFID|temp_imemload_output [2]),
	.temp_imemload_output_3(\IFID|temp_imemload_output [3]),
	.temp_imemload_output_5(\IFID|temp_imemload_output [5]),
	.Equal31(\CONTROLUNIT|Equal3~1_combout ),
	.temp_imemload_output_15(\IFID|temp_imemload_output [15]),
	.temp_imemload_output_14(\IFID|temp_imemload_output [14]),
	.temp_imemload_output_13(\IFID|temp_imemload_output [13]),
	.temp_imemload_output_12(\IFID|temp_imemload_output [12]),
	.temp_imemload_output_11(\IFID|temp_imemload_output [11]),
	.temp_imemload_output_10(\IFID|temp_imemload_output [10]),
	.temp_imemload_output_9(\IFID|temp_imemload_output [9]),
	.temp_imemload_output_8(\IFID|temp_imemload_output [8]),
	.temp_imemload_output_7(\IFID|temp_imemload_output [7]),
	.temp_imemload_output_6(\IFID|temp_imemload_output [6]),
	.temp_imemload_output_1(\IFID|temp_imemload_output [1]),
	.temp_imemload_output_4(\IFID|temp_imemload_output [4]),
	.Equal32(\CONTROLUNIT|Equal3~9_combout ),
	.WideOr8(\CONTROLUNIT|WideOr8~0_combout ),
	.WideOr2(\CONTROLUNIT|WideOr2~0_combout ),
	.WideOr4(\CONTROLUNIT|WideOr4~0_combout ),
	.WideOr7(\CONTROLUNIT|WideOr7~0_combout ),
	.WideOr1(\CONTROLUNIT|WideOr1~0_combout ),
	.WideOr5(\CONTROLUNIT|WideOr5~0_combout ),
	.WideOr6(\CONTROLUNIT|WideOr6~0_combout ),
	.WideOr0(\CONTROLUNIT|WideOr0~0_combout ),
	.halt_out(\CONTROLUNIT|halt_out~0_combout ),
	.halt_out1(\CONTROLUNIT|halt_out~3_combout ),
	.WideOr3(\CONTROLUNIT|WideOr3~0_combout ),
	.WideOr10(\CONTROLUNIT|WideOr10~0_combout ),
	.memtoreg(\CONTROLUNIT|memtoreg~0_combout ),
	.WideOr9(\CONTROLUNIT|WideOr9~0_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

program_count PC(
	.pccount_1(pccount_1),
	.pccount_0(pccount_0),
	.pccount_2(pccount_2),
	.pccount_3(pccount_3),
	.pccount_5(pccount_5),
	.pccount_4(pccount_4),
	.pccount_7(pccount_7),
	.pccount_6(pccount_6),
	.pccount_9(pccount_9),
	.pccount_8(pccount_8),
	.pccount_11(pccount_11),
	.pccount_10(pccount_10),
	.pccount_13(pccount_13),
	.pccount_12(pccount_12),
	.pccount_15(pccount_15),
	.pccount_14(pccount_14),
	.pccount_17(pccount_17),
	.pccount_16(pccount_16),
	.pccount_19(pccount_19),
	.pccount_18(pccount_18),
	.pccount_20(pccount_20),
	.pccount_21(pccount_21),
	.pccount_23(pccount_23),
	.pccount_22(pccount_22),
	.pccount_25(pccount_25),
	.pccount_24(pccount_24),
	.pccount_26(pccount_26),
	.pccount_27(pccount_27),
	.pccount_29(pccount_29),
	.pccount_28(pccount_28),
	.pccount_31(pccount_31),
	.pccount_30(pccount_30),
	.Mux30(\NPCMUX|Mux30~1_combout ),
	.wen(\HAZARDUNIT|pc_wen~2_combout ),
	.Mux31(\NPCMUX|Mux31~2_combout ),
	.Mux29(\NPCMUX|Mux29~1_combout ),
	.Mux28(\NPCMUX|Mux28~1_combout ),
	.Mux26(\NPCMUX|Mux26~1_combout ),
	.Mux27(\NPCMUX|Mux27~1_combout ),
	.Mux24(\NPCMUX|Mux24~1_combout ),
	.Mux25(\NPCMUX|Mux25~1_combout ),
	.Mux22(\NPCMUX|Mux22~1_combout ),
	.Mux23(\NPCMUX|Mux23~1_combout ),
	.Mux20(\NPCMUX|Mux20~1_combout ),
	.Mux21(\NPCMUX|Mux21~1_combout ),
	.Mux18(\NPCMUX|Mux18~1_combout ),
	.Mux19(\NPCMUX|Mux19~1_combout ),
	.Mux16(\NPCMUX|Mux16~1_combout ),
	.Mux17(\NPCMUX|Mux17~1_combout ),
	.Mux14(\NPCMUX|Mux14~1_combout ),
	.Mux15(\NPCMUX|Mux15~1_combout ),
	.Mux12(\NPCMUX|Mux12~1_combout ),
	.Mux13(\NPCMUX|Mux13~1_combout ),
	.Mux11(\NPCMUX|Mux11~1_combout ),
	.Mux10(\NPCMUX|Mux10~1_combout ),
	.Mux8(\NPCMUX|Mux8~1_combout ),
	.Mux9(\NPCMUX|Mux9~1_combout ),
	.Mux6(\NPCMUX|Mux6~1_combout ),
	.Mux7(\NPCMUX|Mux7~1_combout ),
	.Mux5(\NPCMUX|Mux5~1_combout ),
	.Mux4(\NPCMUX|Mux4~1_combout ),
	.Mux2(\NPCMUX|Mux2~1_combout ),
	.Mux3(\NPCMUX|Mux3~3_combout ),
	.Mux0(\NPCMUX|Mux0~1_combout ),
	.Mux1(\NPCMUX|Mux1~1_combout ),
	.CLK(CPUCLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

register_file REGISTER(
	.temp_regwrite(\MEMWB|temp_regwrite~q ),
	.temp_branchDest_1(\MEMWB|temp_branchDest [1]),
	.temp_branchDest_0(\MEMWB|temp_branchDest [0]),
	.temp_branchDest_3(\MEMWB|temp_branchDest [3]),
	.temp_branchDest_2(\MEMWB|temp_branchDest [2]),
	.temp_branchDest_4(\MEMWB|temp_branchDest [4]),
	.Mux30(\MEMTOREG|Mux30~1_combout ),
	.Mux31(\MEMTOREG|Mux31~1_combout ),
	.Mux29(\MEMTOREG|Mux29~1_combout ),
	.Mux27(\MEMTOREG|Mux27~1_combout ),
	.Mux28(\MEMTOREG|Mux28~1_combout ),
	.Mux23(\MEMTOREG|Mux23~1_combout ),
	.Mux24(\MEMTOREG|Mux24~1_combout ),
	.Mux25(\MEMTOREG|Mux25~1_combout ),
	.Mux26(\MEMTOREG|Mux26~1_combout ),
	.Mux15(\MEMTOREG|Mux15~1_combout ),
	.Mux17(\MEMTOREG|Mux17~1_combout ),
	.Mux16(\MEMTOREG|Mux16~1_combout ),
	.Mux18(\MEMTOREG|Mux18~1_combout ),
	.Mux19(\MEMTOREG|Mux19~1_combout ),
	.Mux21(\MEMTOREG|Mux21~1_combout ),
	.Mux20(\MEMTOREG|Mux20~1_combout ),
	.Mux22(\MEMTOREG|Mux22~1_combout ),
	.Mux0(\MEMTOREG|Mux0~1_combout ),
	.Mux1(\MEMTOREG|Mux1~1_combout ),
	.Mux2(\MEMTOREG|Mux2~1_combout ),
	.Mux5(\MEMTOREG|Mux5~1_combout ),
	.Mux6(\MEMTOREG|Mux6~1_combout ),
	.Mux3(\MEMTOREG|Mux3~1_combout ),
	.Mux4(\MEMTOREG|Mux4~1_combout ),
	.Mux14(\MEMTOREG|Mux14~1_combout ),
	.Mux11(\MEMTOREG|Mux11~1_combout ),
	.Mux12(\MEMTOREG|Mux12~1_combout ),
	.Mux13(\MEMTOREG|Mux13~1_combout ),
	.Mux7(\MEMTOREG|Mux7~1_combout ),
	.Mux8(\MEMTOREG|Mux8~1_combout ),
	.Mux9(\MEMTOREG|Mux9~1_combout ),
	.Mux10(\MEMTOREG|Mux10~1_combout ),
	.temp_imemload_output_17(\IFID|temp_imemload_output [17]),
	.temp_imemload_output_16(\IFID|temp_imemload_output [16]),
	.temp_imemload_output_19(\IFID|temp_imemload_output [19]),
	.temp_imemload_output_18(\IFID|temp_imemload_output [18]),
	.temp_imemload_output_22(\IFID|temp_imemload_output [22]),
	.temp_imemload_output_21(\IFID|temp_imemload_output [21]),
	.temp_imemload_output_24(\IFID|temp_imemload_output [24]),
	.temp_imemload_output_23(\IFID|temp_imemload_output [23]),
	.Mux62(\REGISTER|Mux62~9_combout ),
	.Mux621(\REGISTER|Mux62~19_combout ),
	.Mux301(\REGISTER|Mux30~9_combout ),
	.Mux302(\REGISTER|Mux30~19_combout ),
	.Mux63(\REGISTER|Mux63~9_combout ),
	.Mux631(\REGISTER|Mux63~19_combout ),
	.Mux311(\REGISTER|Mux31~9_combout ),
	.Mux312(\REGISTER|Mux31~19_combout ),
	.Mux291(\REGISTER|Mux29~9_combout ),
	.Mux292(\REGISTER|Mux29~19_combout ),
	.Mux271(\REGISTER|Mux27~9_combout ),
	.Mux272(\REGISTER|Mux27~19_combout ),
	.Mux281(\REGISTER|Mux28~9_combout ),
	.Mux282(\REGISTER|Mux28~19_combout ),
	.Mux61(\REGISTER|Mux61~9_combout ),
	.Mux611(\REGISTER|Mux61~19_combout ),
	.Mux231(\REGISTER|Mux23~9_combout ),
	.Mux232(\REGISTER|Mux23~19_combout ),
	.Mux241(\REGISTER|Mux24~9_combout ),
	.Mux242(\REGISTER|Mux24~19_combout ),
	.Mux251(\REGISTER|Mux25~9_combout ),
	.Mux252(\REGISTER|Mux25~19_combout ),
	.Mux261(\REGISTER|Mux26~9_combout ),
	.Mux262(\REGISTER|Mux26~19_combout ),
	.Mux60(\REGISTER|Mux60~9_combout ),
	.Mux601(\REGISTER|Mux60~19_combout ),
	.Mux151(\REGISTER|Mux15~9_combout ),
	.Mux152(\REGISTER|Mux15~19_combout ),
	.Mux171(\REGISTER|Mux17~9_combout ),
	.Mux172(\REGISTER|Mux17~19_combout ),
	.Mux161(\REGISTER|Mux16~9_combout ),
	.Mux162(\REGISTER|Mux16~19_combout ),
	.Mux181(\REGISTER|Mux18~9_combout ),
	.Mux182(\REGISTER|Mux18~19_combout ),
	.Mux191(\REGISTER|Mux19~9_combout ),
	.Mux192(\REGISTER|Mux19~19_combout ),
	.Mux211(\REGISTER|Mux21~9_combout ),
	.Mux212(\REGISTER|Mux21~19_combout ),
	.Mux201(\REGISTER|Mux20~9_combout ),
	.Mux202(\REGISTER|Mux20~19_combout ),
	.Mux221(\REGISTER|Mux22~9_combout ),
	.Mux222(\REGISTER|Mux22~19_combout ),
	.Mux59(\REGISTER|Mux59~9_combout ),
	.Mux591(\REGISTER|Mux59~19_combout ),
	.Mux01(\REGISTER|Mux0~9_combout ),
	.Mux02(\REGISTER|Mux0~19_combout ),
	.Mux110(\REGISTER|Mux1~9_combout ),
	.Mux111(\REGISTER|Mux1~19_combout ),
	.Mux210(\REGISTER|Mux2~9_combout ),
	.Mux213(\REGISTER|Mux2~19_combout ),
	.Mux51(\REGISTER|Mux5~9_combout ),
	.Mux52(\REGISTER|Mux5~19_combout ),
	.Mux64(\REGISTER|Mux6~9_combout ),
	.Mux65(\REGISTER|Mux6~19_combout ),
	.Mux32(\REGISTER|Mux3~9_combout ),
	.Mux33(\REGISTER|Mux3~19_combout ),
	.Mux41(\REGISTER|Mux4~9_combout ),
	.Mux42(\REGISTER|Mux4~19_combout ),
	.Mux141(\REGISTER|Mux14~9_combout ),
	.Mux142(\REGISTER|Mux14~19_combout ),
	.Mux112(\REGISTER|Mux11~9_combout ),
	.Mux113(\REGISTER|Mux11~19_combout ),
	.Mux121(\REGISTER|Mux12~9_combout ),
	.Mux122(\REGISTER|Mux12~19_combout ),
	.Mux131(\REGISTER|Mux13~9_combout ),
	.Mux132(\REGISTER|Mux13~19_combout ),
	.Mux71(\REGISTER|Mux7~9_combout ),
	.Mux72(\REGISTER|Mux7~19_combout ),
	.Mux81(\REGISTER|Mux8~9_combout ),
	.Mux82(\REGISTER|Mux8~19_combout ),
	.Mux91(\REGISTER|Mux9~9_combout ),
	.Mux92(\REGISTER|Mux9~19_combout ),
	.Mux101(\REGISTER|Mux10~9_combout ),
	.Mux102(\REGISTER|Mux10~19_combout ),
	.Mux48(\REGISTER|Mux48~9_combout ),
	.Mux481(\REGISTER|Mux48~19_combout ),
	.Mux511(\REGISTER|Mux51~9_combout ),
	.Mux512(\REGISTER|Mux51~19_combout ),
	.Mux36(\REGISTER|Mux36~9_combout ),
	.Mux361(\REGISTER|Mux36~19_combout ),
	.Mux45(\REGISTER|Mux45~9_combout ),
	.Mux451(\REGISTER|Mux45~19_combout ),
	.Mux46(\REGISTER|Mux46~9_combout ),
	.Mux461(\REGISTER|Mux46~19_combout ),
	.Mux47(\REGISTER|Mux47~9_combout ),
	.Mux471(\REGISTER|Mux47~19_combout ),
	.Mux321(\REGISTER|Mux32~9_combout ),
	.Mux322(\REGISTER|Mux32~19_combout ),
	.Mux331(\REGISTER|Mux33~9_combout ),
	.Mux332(\REGISTER|Mux33~19_combout ),
	.Mux34(\REGISTER|Mux34~9_combout ),
	.Mux341(\REGISTER|Mux34~19_combout ),
	.Mux35(\REGISTER|Mux35~9_combout ),
	.Mux351(\REGISTER|Mux35~19_combout ),
	.Mux37(\REGISTER|Mux37~9_combout ),
	.Mux371(\REGISTER|Mux37~19_combout ),
	.Mux38(\REGISTER|Mux38~9_combout ),
	.Mux381(\REGISTER|Mux38~19_combout ),
	.Mux39(\REGISTER|Mux39~9_combout ),
	.Mux391(\REGISTER|Mux39~19_combout ),
	.Mux40(\REGISTER|Mux40~9_combout ),
	.Mux401(\REGISTER|Mux40~19_combout ),
	.Mux411(\REGISTER|Mux41~9_combout ),
	.Mux412(\REGISTER|Mux41~19_combout ),
	.Mux421(\REGISTER|Mux42~9_combout ),
	.Mux422(\REGISTER|Mux42~19_combout ),
	.Mux43(\REGISTER|Mux43~9_combout ),
	.Mux431(\REGISTER|Mux43~19_combout ),
	.Mux44(\REGISTER|Mux44~9_combout ),
	.Mux441(\REGISTER|Mux44~19_combout ),
	.Mux53(\REGISTER|Mux53~9_combout ),
	.Mux531(\REGISTER|Mux53~19_combout ),
	.Mux49(\REGISTER|Mux49~9_combout ),
	.Mux491(\REGISTER|Mux49~19_combout ),
	.Mux54(\REGISTER|Mux54~9_combout ),
	.Mux541(\REGISTER|Mux54~19_combout ),
	.Mux55(\REGISTER|Mux55~9_combout ),
	.Mux551(\REGISTER|Mux55~19_combout ),
	.Mux56(\REGISTER|Mux56~9_combout ),
	.Mux561(\REGISTER|Mux56~19_combout ),
	.Mux57(\REGISTER|Mux57~9_combout ),
	.Mux571(\REGISTER|Mux57~19_combout ),
	.Mux58(\REGISTER|Mux58~9_combout ),
	.Mux581(\REGISTER|Mux58~19_combout ),
	.Mux50(\REGISTER|Mux50~9_combout ),
	.Mux501(\REGISTER|Mux50~19_combout ),
	.Mux521(\REGISTER|Mux52~9_combout ),
	.Mux522(\REGISTER|Mux52~19_combout ),
	.CLK(CPUCLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X62_Y45_N2
cycloneive_lcell_comb \branch_count_output[2]~0 (
// Equation(s):
// \branch_count_output[2]~0_combout  = (temp_npc_2 & (temp_iMemLoad_0 $ (VCC))) # (!temp_npc_2 & (temp_iMemLoad_0 & VCC))
// \branch_count_output[2]~1  = CARRY((temp_npc_2 & temp_iMemLoad_0))

	.dataa(\EXMEM|temp_npc [2]),
	.datab(\EXMEM|temp_iMemLoad [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\branch_count_output[2]~0_combout ),
	.cout(\branch_count_output[2]~1 ));
// synopsys translate_off
defparam \branch_count_output[2]~0 .lut_mask = 16'h6688;
defparam \branch_count_output[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N2
cycloneive_lcell_comb \pc_count_four_output[2]~0 (
// Equation(s):
// \pc_count_four_output[2]~0_combout  = pccount_2 $ (VCC)
// \pc_count_four_output[2]~1  = CARRY(pccount_2)

	.dataa(pccount_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\pc_count_four_output[2]~0_combout ),
	.cout(\pc_count_four_output[2]~1 ));
// synopsys translate_off
defparam \pc_count_four_output[2]~0 .lut_mask = 16'h55AA;
defparam \pc_count_four_output[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N4
cycloneive_lcell_comb \pc_count_four_output[3]~2 (
// Equation(s):
// \pc_count_four_output[3]~2_combout  = (pccount_3 & (!\pc_count_four_output[2]~1 )) # (!pccount_3 & ((\pc_count_four_output[2]~1 ) # (GND)))
// \pc_count_four_output[3]~3  = CARRY((!\pc_count_four_output[2]~1 ) # (!pccount_3))

	.dataa(pccount_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[2]~1 ),
	.combout(\pc_count_four_output[3]~2_combout ),
	.cout(\pc_count_four_output[3]~3 ));
// synopsys translate_off
defparam \pc_count_four_output[3]~2 .lut_mask = 16'h5A5F;
defparam \pc_count_four_output[3]~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N4
cycloneive_lcell_comb \branch_count_output[3]~2 (
// Equation(s):
// \branch_count_output[3]~2_combout  = (temp_npc_3 & ((temp_iMemLoad_1 & (\branch_count_output[2]~1  & VCC)) # (!temp_iMemLoad_1 & (!\branch_count_output[2]~1 )))) # (!temp_npc_3 & ((temp_iMemLoad_1 & (!\branch_count_output[2]~1 )) # (!temp_iMemLoad_1 & 
// ((\branch_count_output[2]~1 ) # (GND)))))
// \branch_count_output[3]~3  = CARRY((temp_npc_3 & (!temp_iMemLoad_1 & !\branch_count_output[2]~1 )) # (!temp_npc_3 & ((!\branch_count_output[2]~1 ) # (!temp_iMemLoad_1))))

	.dataa(\EXMEM|temp_npc [3]),
	.datab(\EXMEM|temp_iMemLoad [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[2]~1 ),
	.combout(\branch_count_output[3]~2_combout ),
	.cout(\branch_count_output[3]~3 ));
// synopsys translate_off
defparam \branch_count_output[3]~2 .lut_mask = 16'h9617;
defparam \branch_count_output[3]~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N6
cycloneive_lcell_comb \pc_count_four_output[4]~4 (
// Equation(s):
// \pc_count_four_output[4]~4_combout  = (pccount_4 & (\pc_count_four_output[3]~3  $ (GND))) # (!pccount_4 & (!\pc_count_four_output[3]~3  & VCC))
// \pc_count_four_output[4]~5  = CARRY((pccount_4 & !\pc_count_four_output[3]~3 ))

	.dataa(gnd),
	.datab(pccount_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[3]~3 ),
	.combout(\pc_count_four_output[4]~4_combout ),
	.cout(\pc_count_four_output[4]~5 ));
// synopsys translate_off
defparam \pc_count_four_output[4]~4 .lut_mask = 16'hC30C;
defparam \pc_count_four_output[4]~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N8
cycloneive_lcell_comb \pc_count_four_output[5]~6 (
// Equation(s):
// \pc_count_four_output[5]~6_combout  = (pccount_5 & (!\pc_count_four_output[4]~5 )) # (!pccount_5 & ((\pc_count_four_output[4]~5 ) # (GND)))
// \pc_count_four_output[5]~7  = CARRY((!\pc_count_four_output[4]~5 ) # (!pccount_5))

	.dataa(pccount_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[4]~5 ),
	.combout(\pc_count_four_output[5]~6_combout ),
	.cout(\pc_count_four_output[5]~7 ));
// synopsys translate_off
defparam \pc_count_four_output[5]~6 .lut_mask = 16'h5A5F;
defparam \pc_count_four_output[5]~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N6
cycloneive_lcell_comb \branch_count_output[4]~4 (
// Equation(s):
// \branch_count_output[4]~4_combout  = ((temp_iMemLoad_2 $ (temp_npc_4 $ (!\branch_count_output[3]~3 )))) # (GND)
// \branch_count_output[4]~5  = CARRY((temp_iMemLoad_2 & ((temp_npc_4) # (!\branch_count_output[3]~3 ))) # (!temp_iMemLoad_2 & (temp_npc_4 & !\branch_count_output[3]~3 )))

	.dataa(\EXMEM|temp_iMemLoad [2]),
	.datab(\EXMEM|temp_npc [4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[3]~3 ),
	.combout(\branch_count_output[4]~4_combout ),
	.cout(\branch_count_output[4]~5 ));
// synopsys translate_off
defparam \branch_count_output[4]~4 .lut_mask = 16'h698E;
defparam \branch_count_output[4]~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N8
cycloneive_lcell_comb \branch_count_output[5]~6 (
// Equation(s):
// \branch_count_output[5]~6_combout  = (temp_npc_5 & ((temp_iMemLoad_3 & (\branch_count_output[4]~5  & VCC)) # (!temp_iMemLoad_3 & (!\branch_count_output[4]~5 )))) # (!temp_npc_5 & ((temp_iMemLoad_3 & (!\branch_count_output[4]~5 )) # (!temp_iMemLoad_3 & 
// ((\branch_count_output[4]~5 ) # (GND)))))
// \branch_count_output[5]~7  = CARRY((temp_npc_5 & (!temp_iMemLoad_3 & !\branch_count_output[4]~5 )) # (!temp_npc_5 & ((!\branch_count_output[4]~5 ) # (!temp_iMemLoad_3))))

	.dataa(\EXMEM|temp_npc [5]),
	.datab(\EXMEM|temp_iMemLoad [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[4]~5 ),
	.combout(\branch_count_output[5]~6_combout ),
	.cout(\branch_count_output[5]~7 ));
// synopsys translate_off
defparam \branch_count_output[5]~6 .lut_mask = 16'h9617;
defparam \branch_count_output[5]~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N10
cycloneive_lcell_comb \pc_count_four_output[6]~8 (
// Equation(s):
// \pc_count_four_output[6]~8_combout  = (pccount_6 & (\pc_count_four_output[5]~7  $ (GND))) # (!pccount_6 & (!\pc_count_four_output[5]~7  & VCC))
// \pc_count_four_output[6]~9  = CARRY((pccount_6 & !\pc_count_four_output[5]~7 ))

	.dataa(gnd),
	.datab(pccount_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[5]~7 ),
	.combout(\pc_count_four_output[6]~8_combout ),
	.cout(\pc_count_four_output[6]~9 ));
// synopsys translate_off
defparam \pc_count_four_output[6]~8 .lut_mask = 16'hC30C;
defparam \pc_count_four_output[6]~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N12
cycloneive_lcell_comb \pc_count_four_output[7]~10 (
// Equation(s):
// \pc_count_four_output[7]~10_combout  = (pccount_7 & (!\pc_count_four_output[6]~9 )) # (!pccount_7 & ((\pc_count_four_output[6]~9 ) # (GND)))
// \pc_count_four_output[7]~11  = CARRY((!\pc_count_four_output[6]~9 ) # (!pccount_7))

	.dataa(pccount_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[6]~9 ),
	.combout(\pc_count_four_output[7]~10_combout ),
	.cout(\pc_count_four_output[7]~11 ));
// synopsys translate_off
defparam \pc_count_four_output[7]~10 .lut_mask = 16'h5A5F;
defparam \pc_count_four_output[7]~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N10
cycloneive_lcell_comb \branch_count_output[6]~8 (
// Equation(s):
// \branch_count_output[6]~8_combout  = ((temp_npc_6 $ (temp_iMemLoad_4 $ (!\branch_count_output[5]~7 )))) # (GND)
// \branch_count_output[6]~9  = CARRY((temp_npc_6 & ((temp_iMemLoad_4) # (!\branch_count_output[5]~7 ))) # (!temp_npc_6 & (temp_iMemLoad_4 & !\branch_count_output[5]~7 )))

	.dataa(\EXMEM|temp_npc [6]),
	.datab(\EXMEM|temp_iMemLoad [4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[5]~7 ),
	.combout(\branch_count_output[6]~8_combout ),
	.cout(\branch_count_output[6]~9 ));
// synopsys translate_off
defparam \branch_count_output[6]~8 .lut_mask = 16'h698E;
defparam \branch_count_output[6]~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N12
cycloneive_lcell_comb \branch_count_output[7]~10 (
// Equation(s):
// \branch_count_output[7]~10_combout  = (temp_npc_7 & ((temp_iMemLoad_5 & (\branch_count_output[6]~9  & VCC)) # (!temp_iMemLoad_5 & (!\branch_count_output[6]~9 )))) # (!temp_npc_7 & ((temp_iMemLoad_5 & (!\branch_count_output[6]~9 )) # (!temp_iMemLoad_5 & 
// ((\branch_count_output[6]~9 ) # (GND)))))
// \branch_count_output[7]~11  = CARRY((temp_npc_7 & (!temp_iMemLoad_5 & !\branch_count_output[6]~9 )) # (!temp_npc_7 & ((!\branch_count_output[6]~9 ) # (!temp_iMemLoad_5))))

	.dataa(\EXMEM|temp_npc [7]),
	.datab(\EXMEM|temp_iMemLoad [5]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[6]~9 ),
	.combout(\branch_count_output[7]~10_combout ),
	.cout(\branch_count_output[7]~11 ));
// synopsys translate_off
defparam \branch_count_output[7]~10 .lut_mask = 16'h9617;
defparam \branch_count_output[7]~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N14
cycloneive_lcell_comb \pc_count_four_output[8]~12 (
// Equation(s):
// \pc_count_four_output[8]~12_combout  = (pccount_8 & (\pc_count_four_output[7]~11  $ (GND))) # (!pccount_8 & (!\pc_count_four_output[7]~11  & VCC))
// \pc_count_four_output[8]~13  = CARRY((pccount_8 & !\pc_count_four_output[7]~11 ))

	.dataa(pccount_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[7]~11 ),
	.combout(\pc_count_four_output[8]~12_combout ),
	.cout(\pc_count_four_output[8]~13 ));
// synopsys translate_off
defparam \pc_count_four_output[8]~12 .lut_mask = 16'hA50A;
defparam \pc_count_four_output[8]~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N16
cycloneive_lcell_comb \pc_count_four_output[9]~14 (
// Equation(s):
// \pc_count_four_output[9]~14_combout  = (pccount_9 & (!\pc_count_four_output[8]~13 )) # (!pccount_9 & ((\pc_count_four_output[8]~13 ) # (GND)))
// \pc_count_four_output[9]~15  = CARRY((!\pc_count_four_output[8]~13 ) # (!pccount_9))

	.dataa(pccount_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[8]~13 ),
	.combout(\pc_count_four_output[9]~14_combout ),
	.cout(\pc_count_four_output[9]~15 ));
// synopsys translate_off
defparam \pc_count_four_output[9]~14 .lut_mask = 16'h5A5F;
defparam \pc_count_four_output[9]~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N14
cycloneive_lcell_comb \branch_count_output[8]~12 (
// Equation(s):
// \branch_count_output[8]~12_combout  = ((temp_iMemLoad_6 $ (temp_npc_8 $ (!\branch_count_output[7]~11 )))) # (GND)
// \branch_count_output[8]~13  = CARRY((temp_iMemLoad_6 & ((temp_npc_8) # (!\branch_count_output[7]~11 ))) # (!temp_iMemLoad_6 & (temp_npc_8 & !\branch_count_output[7]~11 )))

	.dataa(\EXMEM|temp_iMemLoad [6]),
	.datab(\EXMEM|temp_npc [8]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[7]~11 ),
	.combout(\branch_count_output[8]~12_combout ),
	.cout(\branch_count_output[8]~13 ));
// synopsys translate_off
defparam \branch_count_output[8]~12 .lut_mask = 16'h698E;
defparam \branch_count_output[8]~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N16
cycloneive_lcell_comb \branch_count_output[9]~14 (
// Equation(s):
// \branch_count_output[9]~14_combout  = (temp_npc_9 & ((temp_iMemLoad_7 & (\branch_count_output[8]~13  & VCC)) # (!temp_iMemLoad_7 & (!\branch_count_output[8]~13 )))) # (!temp_npc_9 & ((temp_iMemLoad_7 & (!\branch_count_output[8]~13 )) # (!temp_iMemLoad_7 & 
// ((\branch_count_output[8]~13 ) # (GND)))))
// \branch_count_output[9]~15  = CARRY((temp_npc_9 & (!temp_iMemLoad_7 & !\branch_count_output[8]~13 )) # (!temp_npc_9 & ((!\branch_count_output[8]~13 ) # (!temp_iMemLoad_7))))

	.dataa(\EXMEM|temp_npc [9]),
	.datab(\EXMEM|temp_iMemLoad [7]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[8]~13 ),
	.combout(\branch_count_output[9]~14_combout ),
	.cout(\branch_count_output[9]~15 ));
// synopsys translate_off
defparam \branch_count_output[9]~14 .lut_mask = 16'h9617;
defparam \branch_count_output[9]~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N18
cycloneive_lcell_comb \pc_count_four_output[10]~16 (
// Equation(s):
// \pc_count_four_output[10]~16_combout  = (pccount_10 & (\pc_count_four_output[9]~15  $ (GND))) # (!pccount_10 & (!\pc_count_four_output[9]~15  & VCC))
// \pc_count_four_output[10]~17  = CARRY((pccount_10 & !\pc_count_four_output[9]~15 ))

	.dataa(pccount_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[9]~15 ),
	.combout(\pc_count_four_output[10]~16_combout ),
	.cout(\pc_count_four_output[10]~17 ));
// synopsys translate_off
defparam \pc_count_four_output[10]~16 .lut_mask = 16'hA50A;
defparam \pc_count_four_output[10]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N20
cycloneive_lcell_comb \pc_count_four_output[11]~18 (
// Equation(s):
// \pc_count_four_output[11]~18_combout  = (pccount_11 & (!\pc_count_four_output[10]~17 )) # (!pccount_11 & ((\pc_count_four_output[10]~17 ) # (GND)))
// \pc_count_four_output[11]~19  = CARRY((!\pc_count_four_output[10]~17 ) # (!pccount_11))

	.dataa(gnd),
	.datab(pccount_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[10]~17 ),
	.combout(\pc_count_four_output[11]~18_combout ),
	.cout(\pc_count_four_output[11]~19 ));
// synopsys translate_off
defparam \pc_count_four_output[11]~18 .lut_mask = 16'h3C3F;
defparam \pc_count_four_output[11]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N18
cycloneive_lcell_comb \branch_count_output[10]~16 (
// Equation(s):
// \branch_count_output[10]~16_combout  = ((temp_npc_10 $ (temp_iMemLoad_8 $ (!\branch_count_output[9]~15 )))) # (GND)
// \branch_count_output[10]~17  = CARRY((temp_npc_10 & ((temp_iMemLoad_8) # (!\branch_count_output[9]~15 ))) # (!temp_npc_10 & (temp_iMemLoad_8 & !\branch_count_output[9]~15 )))

	.dataa(\EXMEM|temp_npc [10]),
	.datab(\EXMEM|temp_iMemLoad [8]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[9]~15 ),
	.combout(\branch_count_output[10]~16_combout ),
	.cout(\branch_count_output[10]~17 ));
// synopsys translate_off
defparam \branch_count_output[10]~16 .lut_mask = 16'h698E;
defparam \branch_count_output[10]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N20
cycloneive_lcell_comb \branch_count_output[11]~18 (
// Equation(s):
// \branch_count_output[11]~18_combout  = (temp_iMemLoad_9 & ((temp_npc_11 & (\branch_count_output[10]~17  & VCC)) # (!temp_npc_11 & (!\branch_count_output[10]~17 )))) # (!temp_iMemLoad_9 & ((temp_npc_11 & (!\branch_count_output[10]~17 )) # (!temp_npc_11 & 
// ((\branch_count_output[10]~17 ) # (GND)))))
// \branch_count_output[11]~19  = CARRY((temp_iMemLoad_9 & (!temp_npc_11 & !\branch_count_output[10]~17 )) # (!temp_iMemLoad_9 & ((!\branch_count_output[10]~17 ) # (!temp_npc_11))))

	.dataa(\EXMEM|temp_iMemLoad [9]),
	.datab(\EXMEM|temp_npc [11]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[10]~17 ),
	.combout(\branch_count_output[11]~18_combout ),
	.cout(\branch_count_output[11]~19 ));
// synopsys translate_off
defparam \branch_count_output[11]~18 .lut_mask = 16'h9617;
defparam \branch_count_output[11]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N22
cycloneive_lcell_comb \pc_count_four_output[12]~20 (
// Equation(s):
// \pc_count_four_output[12]~20_combout  = (pccount_12 & (\pc_count_four_output[11]~19  $ (GND))) # (!pccount_12 & (!\pc_count_four_output[11]~19  & VCC))
// \pc_count_four_output[12]~21  = CARRY((pccount_12 & !\pc_count_four_output[11]~19 ))

	.dataa(pccount_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[11]~19 ),
	.combout(\pc_count_four_output[12]~20_combout ),
	.cout(\pc_count_four_output[12]~21 ));
// synopsys translate_off
defparam \pc_count_four_output[12]~20 .lut_mask = 16'hA50A;
defparam \pc_count_four_output[12]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N24
cycloneive_lcell_comb \pc_count_four_output[13]~22 (
// Equation(s):
// \pc_count_four_output[13]~22_combout  = (pccount_13 & (!\pc_count_four_output[12]~21 )) # (!pccount_13 & ((\pc_count_four_output[12]~21 ) # (GND)))
// \pc_count_four_output[13]~23  = CARRY((!\pc_count_four_output[12]~21 ) # (!pccount_13))

	.dataa(pccount_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[12]~21 ),
	.combout(\pc_count_four_output[13]~22_combout ),
	.cout(\pc_count_four_output[13]~23 ));
// synopsys translate_off
defparam \pc_count_four_output[13]~22 .lut_mask = 16'h5A5F;
defparam \pc_count_four_output[13]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N22
cycloneive_lcell_comb \branch_count_output[12]~20 (
// Equation(s):
// \branch_count_output[12]~20_combout  = ((temp_iMemLoad_10 $ (temp_npc_12 $ (!\branch_count_output[11]~19 )))) # (GND)
// \branch_count_output[12]~21  = CARRY((temp_iMemLoad_10 & ((temp_npc_12) # (!\branch_count_output[11]~19 ))) # (!temp_iMemLoad_10 & (temp_npc_12 & !\branch_count_output[11]~19 )))

	.dataa(\EXMEM|temp_iMemLoad [10]),
	.datab(\EXMEM|temp_npc [12]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[11]~19 ),
	.combout(\branch_count_output[12]~20_combout ),
	.cout(\branch_count_output[12]~21 ));
// synopsys translate_off
defparam \branch_count_output[12]~20 .lut_mask = 16'h698E;
defparam \branch_count_output[12]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N24
cycloneive_lcell_comb \branch_count_output[13]~22 (
// Equation(s):
// \branch_count_output[13]~22_combout  = (temp_npc_13 & ((temp_iMemLoad_11 & (\branch_count_output[12]~21  & VCC)) # (!temp_iMemLoad_11 & (!\branch_count_output[12]~21 )))) # (!temp_npc_13 & ((temp_iMemLoad_11 & (!\branch_count_output[12]~21 )) # 
// (!temp_iMemLoad_11 & ((\branch_count_output[12]~21 ) # (GND)))))
// \branch_count_output[13]~23  = CARRY((temp_npc_13 & (!temp_iMemLoad_11 & !\branch_count_output[12]~21 )) # (!temp_npc_13 & ((!\branch_count_output[12]~21 ) # (!temp_iMemLoad_11))))

	.dataa(\EXMEM|temp_npc [13]),
	.datab(\EXMEM|temp_iMemLoad [11]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[12]~21 ),
	.combout(\branch_count_output[13]~22_combout ),
	.cout(\branch_count_output[13]~23 ));
// synopsys translate_off
defparam \branch_count_output[13]~22 .lut_mask = 16'h9617;
defparam \branch_count_output[13]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N26
cycloneive_lcell_comb \pc_count_four_output[14]~24 (
// Equation(s):
// \pc_count_four_output[14]~24_combout  = (pccount_14 & (\pc_count_four_output[13]~23  $ (GND))) # (!pccount_14 & (!\pc_count_four_output[13]~23  & VCC))
// \pc_count_four_output[14]~25  = CARRY((pccount_14 & !\pc_count_four_output[13]~23 ))

	.dataa(gnd),
	.datab(pccount_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[13]~23 ),
	.combout(\pc_count_four_output[14]~24_combout ),
	.cout(\pc_count_four_output[14]~25 ));
// synopsys translate_off
defparam \pc_count_four_output[14]~24 .lut_mask = 16'hC30C;
defparam \pc_count_four_output[14]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N28
cycloneive_lcell_comb \pc_count_four_output[15]~26 (
// Equation(s):
// \pc_count_four_output[15]~26_combout  = (pccount_15 & (!\pc_count_four_output[14]~25 )) # (!pccount_15 & ((\pc_count_four_output[14]~25 ) # (GND)))
// \pc_count_four_output[15]~27  = CARRY((!\pc_count_four_output[14]~25 ) # (!pccount_15))

	.dataa(gnd),
	.datab(pccount_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[14]~25 ),
	.combout(\pc_count_four_output[15]~26_combout ),
	.cout(\pc_count_four_output[15]~27 ));
// synopsys translate_off
defparam \pc_count_four_output[15]~26 .lut_mask = 16'h3C3F;
defparam \pc_count_four_output[15]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N26
cycloneive_lcell_comb \branch_count_output[14]~24 (
// Equation(s):
// \branch_count_output[14]~24_combout  = ((temp_iMemLoad_12 $ (temp_npc_14 $ (!\branch_count_output[13]~23 )))) # (GND)
// \branch_count_output[14]~25  = CARRY((temp_iMemLoad_12 & ((temp_npc_14) # (!\branch_count_output[13]~23 ))) # (!temp_iMemLoad_12 & (temp_npc_14 & !\branch_count_output[13]~23 )))

	.dataa(\EXMEM|temp_iMemLoad [12]),
	.datab(\EXMEM|temp_npc [14]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[13]~23 ),
	.combout(\branch_count_output[14]~24_combout ),
	.cout(\branch_count_output[14]~25 ));
// synopsys translate_off
defparam \branch_count_output[14]~24 .lut_mask = 16'h698E;
defparam \branch_count_output[14]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N28
cycloneive_lcell_comb \branch_count_output[15]~26 (
// Equation(s):
// \branch_count_output[15]~26_combout  = (temp_iMemLoad_13 & ((temp_npc_15 & (\branch_count_output[14]~25  & VCC)) # (!temp_npc_15 & (!\branch_count_output[14]~25 )))) # (!temp_iMemLoad_13 & ((temp_npc_15 & (!\branch_count_output[14]~25 )) # (!temp_npc_15 & 
// ((\branch_count_output[14]~25 ) # (GND)))))
// \branch_count_output[15]~27  = CARRY((temp_iMemLoad_13 & (!temp_npc_15 & !\branch_count_output[14]~25 )) # (!temp_iMemLoad_13 & ((!\branch_count_output[14]~25 ) # (!temp_npc_15))))

	.dataa(\EXMEM|temp_iMemLoad [13]),
	.datab(\EXMEM|temp_npc [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[14]~25 ),
	.combout(\branch_count_output[15]~26_combout ),
	.cout(\branch_count_output[15]~27 ));
// synopsys translate_off
defparam \branch_count_output[15]~26 .lut_mask = 16'h9617;
defparam \branch_count_output[15]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N30
cycloneive_lcell_comb \pc_count_four_output[16]~28 (
// Equation(s):
// \pc_count_four_output[16]~28_combout  = (pccount_16 & (\pc_count_four_output[15]~27  $ (GND))) # (!pccount_16 & (!\pc_count_four_output[15]~27  & VCC))
// \pc_count_four_output[16]~29  = CARRY((pccount_16 & !\pc_count_four_output[15]~27 ))

	.dataa(gnd),
	.datab(pccount_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[15]~27 ),
	.combout(\pc_count_four_output[16]~28_combout ),
	.cout(\pc_count_four_output[16]~29 ));
// synopsys translate_off
defparam \pc_count_four_output[16]~28 .lut_mask = 16'hC30C;
defparam \pc_count_four_output[16]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N0
cycloneive_lcell_comb \pc_count_four_output[17]~30 (
// Equation(s):
// \pc_count_four_output[17]~30_combout  = (pccount_17 & (!\pc_count_four_output[16]~29 )) # (!pccount_17 & ((\pc_count_four_output[16]~29 ) # (GND)))
// \pc_count_four_output[17]~31  = CARRY((!\pc_count_four_output[16]~29 ) # (!pccount_17))

	.dataa(gnd),
	.datab(pccount_17),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[16]~29 ),
	.combout(\pc_count_four_output[17]~30_combout ),
	.cout(\pc_count_four_output[17]~31 ));
// synopsys translate_off
defparam \pc_count_four_output[17]~30 .lut_mask = 16'h3C3F;
defparam \pc_count_four_output[17]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N30
cycloneive_lcell_comb \branch_count_output[16]~28 (
// Equation(s):
// \branch_count_output[16]~28_combout  = ((temp_npc_16 $ (temp_iMemLoad_14 $ (!\branch_count_output[15]~27 )))) # (GND)
// \branch_count_output[16]~29  = CARRY((temp_npc_16 & ((temp_iMemLoad_14) # (!\branch_count_output[15]~27 ))) # (!temp_npc_16 & (temp_iMemLoad_14 & !\branch_count_output[15]~27 )))

	.dataa(\EXMEM|temp_npc [16]),
	.datab(\EXMEM|temp_iMemLoad [14]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[15]~27 ),
	.combout(\branch_count_output[16]~28_combout ),
	.cout(\branch_count_output[16]~29 ));
// synopsys translate_off
defparam \branch_count_output[16]~28 .lut_mask = 16'h698E;
defparam \branch_count_output[16]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N0
cycloneive_lcell_comb \branch_count_output[17]~30 (
// Equation(s):
// \branch_count_output[17]~30_combout  = (temp_iMemLoad_15 & ((temp_npc_17 & (\branch_count_output[16]~29  & VCC)) # (!temp_npc_17 & (!\branch_count_output[16]~29 )))) # (!temp_iMemLoad_15 & ((temp_npc_17 & (!\branch_count_output[16]~29 )) # (!temp_npc_17 & 
// ((\branch_count_output[16]~29 ) # (GND)))))
// \branch_count_output[17]~31  = CARRY((temp_iMemLoad_15 & (!temp_npc_17 & !\branch_count_output[16]~29 )) # (!temp_iMemLoad_15 & ((!\branch_count_output[16]~29 ) # (!temp_npc_17))))

	.dataa(\EXMEM|temp_iMemLoad [15]),
	.datab(\EXMEM|temp_npc [17]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[16]~29 ),
	.combout(\branch_count_output[17]~30_combout ),
	.cout(\branch_count_output[17]~31 ));
// synopsys translate_off
defparam \branch_count_output[17]~30 .lut_mask = 16'h9617;
defparam \branch_count_output[17]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N2
cycloneive_lcell_comb \pc_count_four_output[18]~32 (
// Equation(s):
// \pc_count_four_output[18]~32_combout  = (pccount_18 & (\pc_count_four_output[17]~31  $ (GND))) # (!pccount_18 & (!\pc_count_four_output[17]~31  & VCC))
// \pc_count_four_output[18]~33  = CARRY((pccount_18 & !\pc_count_four_output[17]~31 ))

	.dataa(pccount_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[17]~31 ),
	.combout(\pc_count_four_output[18]~32_combout ),
	.cout(\pc_count_four_output[18]~33 ));
// synopsys translate_off
defparam \pc_count_four_output[18]~32 .lut_mask = 16'hA50A;
defparam \pc_count_four_output[18]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N4
cycloneive_lcell_comb \pc_count_four_output[19]~34 (
// Equation(s):
// \pc_count_four_output[19]~34_combout  = (pccount_19 & (!\pc_count_four_output[18]~33 )) # (!pccount_19 & ((\pc_count_four_output[18]~33 ) # (GND)))
// \pc_count_four_output[19]~35  = CARRY((!\pc_count_four_output[18]~33 ) # (!pccount_19))

	.dataa(pccount_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[18]~33 ),
	.combout(\pc_count_four_output[19]~34_combout ),
	.cout(\pc_count_four_output[19]~35 ));
// synopsys translate_off
defparam \pc_count_four_output[19]~34 .lut_mask = 16'h5A5F;
defparam \pc_count_four_output[19]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N2
cycloneive_lcell_comb \branch_count_output[18]~32 (
// Equation(s):
// \branch_count_output[18]~32_combout  = ((temp_signZero_16 $ (temp_npc_18 $ (!\branch_count_output[17]~31 )))) # (GND)
// \branch_count_output[18]~33  = CARRY((temp_signZero_16 & ((temp_npc_18) # (!\branch_count_output[17]~31 ))) # (!temp_signZero_16 & (temp_npc_18 & !\branch_count_output[17]~31 )))

	.dataa(\EXMEM|temp_signZero [16]),
	.datab(\EXMEM|temp_npc [18]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[17]~31 ),
	.combout(\branch_count_output[18]~32_combout ),
	.cout(\branch_count_output[18]~33 ));
// synopsys translate_off
defparam \branch_count_output[18]~32 .lut_mask = 16'h698E;
defparam \branch_count_output[18]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N4
cycloneive_lcell_comb \branch_count_output[19]~34 (
// Equation(s):
// \branch_count_output[19]~34_combout  = (temp_signZero_16 & ((temp_npc_19 & (\branch_count_output[18]~33  & VCC)) # (!temp_npc_19 & (!\branch_count_output[18]~33 )))) # (!temp_signZero_16 & ((temp_npc_19 & (!\branch_count_output[18]~33 )) # (!temp_npc_19 & 
// ((\branch_count_output[18]~33 ) # (GND)))))
// \branch_count_output[19]~35  = CARRY((temp_signZero_16 & (!temp_npc_19 & !\branch_count_output[18]~33 )) # (!temp_signZero_16 & ((!\branch_count_output[18]~33 ) # (!temp_npc_19))))

	.dataa(\EXMEM|temp_signZero [16]),
	.datab(\EXMEM|temp_npc [19]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[18]~33 ),
	.combout(\branch_count_output[19]~34_combout ),
	.cout(\branch_count_output[19]~35 ));
// synopsys translate_off
defparam \branch_count_output[19]~34 .lut_mask = 16'h9617;
defparam \branch_count_output[19]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N6
cycloneive_lcell_comb \branch_count_output[20]~36 (
// Equation(s):
// \branch_count_output[20]~36_combout  = ((temp_signZero_16 $ (temp_npc_20 $ (!\branch_count_output[19]~35 )))) # (GND)
// \branch_count_output[20]~37  = CARRY((temp_signZero_16 & ((temp_npc_20) # (!\branch_count_output[19]~35 ))) # (!temp_signZero_16 & (temp_npc_20 & !\branch_count_output[19]~35 )))

	.dataa(\EXMEM|temp_signZero [16]),
	.datab(\EXMEM|temp_npc [20]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[19]~35 ),
	.combout(\branch_count_output[20]~36_combout ),
	.cout(\branch_count_output[20]~37 ));
// synopsys translate_off
defparam \branch_count_output[20]~36 .lut_mask = 16'h698E;
defparam \branch_count_output[20]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N6
cycloneive_lcell_comb \pc_count_four_output[20]~36 (
// Equation(s):
// \pc_count_four_output[20]~36_combout  = (pccount_20 & (\pc_count_four_output[19]~35  $ (GND))) # (!pccount_20 & (!\pc_count_four_output[19]~35  & VCC))
// \pc_count_four_output[20]~37  = CARRY((pccount_20 & !\pc_count_four_output[19]~35 ))

	.dataa(pccount_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[19]~35 ),
	.combout(\pc_count_four_output[20]~36_combout ),
	.cout(\pc_count_four_output[20]~37 ));
// synopsys translate_off
defparam \pc_count_four_output[20]~36 .lut_mask = 16'hA50A;
defparam \pc_count_four_output[20]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N8
cycloneive_lcell_comb \pc_count_four_output[21]~38 (
// Equation(s):
// \pc_count_four_output[21]~38_combout  = (pccount_21 & (!\pc_count_four_output[20]~37 )) # (!pccount_21 & ((\pc_count_four_output[20]~37 ) # (GND)))
// \pc_count_four_output[21]~39  = CARRY((!\pc_count_four_output[20]~37 ) # (!pccount_21))

	.dataa(gnd),
	.datab(pccount_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[20]~37 ),
	.combout(\pc_count_four_output[21]~38_combout ),
	.cout(\pc_count_four_output[21]~39 ));
// synopsys translate_off
defparam \pc_count_four_output[21]~38 .lut_mask = 16'h3C3F;
defparam \pc_count_four_output[21]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N8
cycloneive_lcell_comb \branch_count_output[21]~38 (
// Equation(s):
// \branch_count_output[21]~38_combout  = (temp_signZero_16 & ((temp_npc_21 & (\branch_count_output[20]~37  & VCC)) # (!temp_npc_21 & (!\branch_count_output[20]~37 )))) # (!temp_signZero_16 & ((temp_npc_21 & (!\branch_count_output[20]~37 )) # (!temp_npc_21 & 
// ((\branch_count_output[20]~37 ) # (GND)))))
// \branch_count_output[21]~39  = CARRY((temp_signZero_16 & (!temp_npc_21 & !\branch_count_output[20]~37 )) # (!temp_signZero_16 & ((!\branch_count_output[20]~37 ) # (!temp_npc_21))))

	.dataa(\EXMEM|temp_signZero [16]),
	.datab(\EXMEM|temp_npc [21]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[20]~37 ),
	.combout(\branch_count_output[21]~38_combout ),
	.cout(\branch_count_output[21]~39 ));
// synopsys translate_off
defparam \branch_count_output[21]~38 .lut_mask = 16'h9617;
defparam \branch_count_output[21]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N10
cycloneive_lcell_comb \pc_count_four_output[22]~40 (
// Equation(s):
// \pc_count_four_output[22]~40_combout  = (pccount_22 & (\pc_count_four_output[21]~39  $ (GND))) # (!pccount_22 & (!\pc_count_four_output[21]~39  & VCC))
// \pc_count_four_output[22]~41  = CARRY((pccount_22 & !\pc_count_four_output[21]~39 ))

	.dataa(pccount_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[21]~39 ),
	.combout(\pc_count_four_output[22]~40_combout ),
	.cout(\pc_count_four_output[22]~41 ));
// synopsys translate_off
defparam \pc_count_four_output[22]~40 .lut_mask = 16'hA50A;
defparam \pc_count_four_output[22]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N12
cycloneive_lcell_comb \pc_count_four_output[23]~42 (
// Equation(s):
// \pc_count_four_output[23]~42_combout  = (pccount_23 & (!\pc_count_four_output[22]~41 )) # (!pccount_23 & ((\pc_count_four_output[22]~41 ) # (GND)))
// \pc_count_four_output[23]~43  = CARRY((!\pc_count_four_output[22]~41 ) # (!pccount_23))

	.dataa(gnd),
	.datab(pccount_23),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[22]~41 ),
	.combout(\pc_count_four_output[23]~42_combout ),
	.cout(\pc_count_four_output[23]~43 ));
// synopsys translate_off
defparam \pc_count_four_output[23]~42 .lut_mask = 16'h3C3F;
defparam \pc_count_four_output[23]~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N10
cycloneive_lcell_comb \branch_count_output[22]~40 (
// Equation(s):
// \branch_count_output[22]~40_combout  = ((temp_signZero_16 $ (temp_npc_22 $ (!\branch_count_output[21]~39 )))) # (GND)
// \branch_count_output[22]~41  = CARRY((temp_signZero_16 & ((temp_npc_22) # (!\branch_count_output[21]~39 ))) # (!temp_signZero_16 & (temp_npc_22 & !\branch_count_output[21]~39 )))

	.dataa(\EXMEM|temp_signZero [16]),
	.datab(\EXMEM|temp_npc [22]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[21]~39 ),
	.combout(\branch_count_output[22]~40_combout ),
	.cout(\branch_count_output[22]~41 ));
// synopsys translate_off
defparam \branch_count_output[22]~40 .lut_mask = 16'h698E;
defparam \branch_count_output[22]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N12
cycloneive_lcell_comb \branch_count_output[23]~42 (
// Equation(s):
// \branch_count_output[23]~42_combout  = (temp_signZero_16 & ((temp_npc_23 & (\branch_count_output[22]~41  & VCC)) # (!temp_npc_23 & (!\branch_count_output[22]~41 )))) # (!temp_signZero_16 & ((temp_npc_23 & (!\branch_count_output[22]~41 )) # (!temp_npc_23 & 
// ((\branch_count_output[22]~41 ) # (GND)))))
// \branch_count_output[23]~43  = CARRY((temp_signZero_16 & (!temp_npc_23 & !\branch_count_output[22]~41 )) # (!temp_signZero_16 & ((!\branch_count_output[22]~41 ) # (!temp_npc_23))))

	.dataa(\EXMEM|temp_signZero [16]),
	.datab(\EXMEM|temp_npc [23]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[22]~41 ),
	.combout(\branch_count_output[23]~42_combout ),
	.cout(\branch_count_output[23]~43 ));
// synopsys translate_off
defparam \branch_count_output[23]~42 .lut_mask = 16'h9617;
defparam \branch_count_output[23]~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N14
cycloneive_lcell_comb \pc_count_four_output[24]~44 (
// Equation(s):
// \pc_count_four_output[24]~44_combout  = (pccount_24 & (\pc_count_four_output[23]~43  $ (GND))) # (!pccount_24 & (!\pc_count_four_output[23]~43  & VCC))
// \pc_count_four_output[24]~45  = CARRY((pccount_24 & !\pc_count_four_output[23]~43 ))

	.dataa(pccount_24),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[23]~43 ),
	.combout(\pc_count_four_output[24]~44_combout ),
	.cout(\pc_count_four_output[24]~45 ));
// synopsys translate_off
defparam \pc_count_four_output[24]~44 .lut_mask = 16'hA50A;
defparam \pc_count_four_output[24]~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N16
cycloneive_lcell_comb \pc_count_four_output[25]~46 (
// Equation(s):
// \pc_count_four_output[25]~46_combout  = (pccount_25 & (!\pc_count_four_output[24]~45 )) # (!pccount_25 & ((\pc_count_four_output[24]~45 ) # (GND)))
// \pc_count_four_output[25]~47  = CARRY((!\pc_count_four_output[24]~45 ) # (!pccount_25))

	.dataa(gnd),
	.datab(pccount_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[24]~45 ),
	.combout(\pc_count_four_output[25]~46_combout ),
	.cout(\pc_count_four_output[25]~47 ));
// synopsys translate_off
defparam \pc_count_four_output[25]~46 .lut_mask = 16'h3C3F;
defparam \pc_count_four_output[25]~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N14
cycloneive_lcell_comb \branch_count_output[24]~44 (
// Equation(s):
// \branch_count_output[24]~44_combout  = ((temp_signZero_16 $ (temp_npc_24 $ (!\branch_count_output[23]~43 )))) # (GND)
// \branch_count_output[24]~45  = CARRY((temp_signZero_16 & ((temp_npc_24) # (!\branch_count_output[23]~43 ))) # (!temp_signZero_16 & (temp_npc_24 & !\branch_count_output[23]~43 )))

	.dataa(\EXMEM|temp_signZero [16]),
	.datab(\EXMEM|temp_npc [24]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[23]~43 ),
	.combout(\branch_count_output[24]~44_combout ),
	.cout(\branch_count_output[24]~45 ));
// synopsys translate_off
defparam \branch_count_output[24]~44 .lut_mask = 16'h698E;
defparam \branch_count_output[24]~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N16
cycloneive_lcell_comb \branch_count_output[25]~46 (
// Equation(s):
// \branch_count_output[25]~46_combout  = (temp_npc_25 & ((temp_signZero_16 & (\branch_count_output[24]~45  & VCC)) # (!temp_signZero_16 & (!\branch_count_output[24]~45 )))) # (!temp_npc_25 & ((temp_signZero_16 & (!\branch_count_output[24]~45 )) # 
// (!temp_signZero_16 & ((\branch_count_output[24]~45 ) # (GND)))))
// \branch_count_output[25]~47  = CARRY((temp_npc_25 & (!temp_signZero_16 & !\branch_count_output[24]~45 )) # (!temp_npc_25 & ((!\branch_count_output[24]~45 ) # (!temp_signZero_16))))

	.dataa(\EXMEM|temp_npc [25]),
	.datab(\EXMEM|temp_signZero [16]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[24]~45 ),
	.combout(\branch_count_output[25]~46_combout ),
	.cout(\branch_count_output[25]~47 ));
// synopsys translate_off
defparam \branch_count_output[25]~46 .lut_mask = 16'h9617;
defparam \branch_count_output[25]~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N18
cycloneive_lcell_comb \branch_count_output[26]~48 (
// Equation(s):
// \branch_count_output[26]~48_combout  = ((temp_npc_26 $ (temp_signZero_16 $ (!\branch_count_output[25]~47 )))) # (GND)
// \branch_count_output[26]~49  = CARRY((temp_npc_26 & ((temp_signZero_16) # (!\branch_count_output[25]~47 ))) # (!temp_npc_26 & (temp_signZero_16 & !\branch_count_output[25]~47 )))

	.dataa(\EXMEM|temp_npc [26]),
	.datab(\EXMEM|temp_signZero [16]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[25]~47 ),
	.combout(\branch_count_output[26]~48_combout ),
	.cout(\branch_count_output[26]~49 ));
// synopsys translate_off
defparam \branch_count_output[26]~48 .lut_mask = 16'h698E;
defparam \branch_count_output[26]~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N18
cycloneive_lcell_comb \pc_count_four_output[26]~48 (
// Equation(s):
// \pc_count_four_output[26]~48_combout  = (pccount_26 & (\pc_count_four_output[25]~47  $ (GND))) # (!pccount_26 & (!\pc_count_four_output[25]~47  & VCC))
// \pc_count_four_output[26]~49  = CARRY((pccount_26 & !\pc_count_four_output[25]~47 ))

	.dataa(pccount_26),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[25]~47 ),
	.combout(\pc_count_four_output[26]~48_combout ),
	.cout(\pc_count_four_output[26]~49 ));
// synopsys translate_off
defparam \pc_count_four_output[26]~48 .lut_mask = 16'hA50A;
defparam \pc_count_four_output[26]~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N20
cycloneive_lcell_comb \pc_count_four_output[27]~50 (
// Equation(s):
// \pc_count_four_output[27]~50_combout  = (pccount_27 & (!\pc_count_four_output[26]~49 )) # (!pccount_27 & ((\pc_count_four_output[26]~49 ) # (GND)))
// \pc_count_four_output[27]~51  = CARRY((!\pc_count_four_output[26]~49 ) # (!pccount_27))

	.dataa(gnd),
	.datab(pccount_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[26]~49 ),
	.combout(\pc_count_four_output[27]~50_combout ),
	.cout(\pc_count_four_output[27]~51 ));
// synopsys translate_off
defparam \pc_count_four_output[27]~50 .lut_mask = 16'h3C3F;
defparam \pc_count_four_output[27]~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N22
cycloneive_lcell_comb \pc_count_four_output[28]~52 (
// Equation(s):
// \pc_count_four_output[28]~52_combout  = (pccount_28 & (\pc_count_four_output[27]~51  $ (GND))) # (!pccount_28 & (!\pc_count_four_output[27]~51  & VCC))
// \pc_count_four_output[28]~53  = CARRY((pccount_28 & !\pc_count_four_output[27]~51 ))

	.dataa(pccount_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[27]~51 ),
	.combout(\pc_count_four_output[28]~52_combout ),
	.cout(\pc_count_four_output[28]~53 ));
// synopsys translate_off
defparam \pc_count_four_output[28]~52 .lut_mask = 16'hA50A;
defparam \pc_count_four_output[28]~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N20
cycloneive_lcell_comb \branch_count_output[27]~50 (
// Equation(s):
// \branch_count_output[27]~50_combout  = (temp_npc_27 & ((temp_signZero_16 & (\branch_count_output[26]~49  & VCC)) # (!temp_signZero_16 & (!\branch_count_output[26]~49 )))) # (!temp_npc_27 & ((temp_signZero_16 & (!\branch_count_output[26]~49 )) # 
// (!temp_signZero_16 & ((\branch_count_output[26]~49 ) # (GND)))))
// \branch_count_output[27]~51  = CARRY((temp_npc_27 & (!temp_signZero_16 & !\branch_count_output[26]~49 )) # (!temp_npc_27 & ((!\branch_count_output[26]~49 ) # (!temp_signZero_16))))

	.dataa(\EXMEM|temp_npc [27]),
	.datab(\EXMEM|temp_signZero [16]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[26]~49 ),
	.combout(\branch_count_output[27]~50_combout ),
	.cout(\branch_count_output[27]~51 ));
// synopsys translate_off
defparam \branch_count_output[27]~50 .lut_mask = 16'h9617;
defparam \branch_count_output[27]~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N24
cycloneive_lcell_comb \pc_count_four_output[29]~54 (
// Equation(s):
// \pc_count_four_output[29]~54_combout  = (pccount_29 & (!\pc_count_four_output[28]~53 )) # (!pccount_29 & ((\pc_count_four_output[28]~53 ) # (GND)))
// \pc_count_four_output[29]~55  = CARRY((!\pc_count_four_output[28]~53 ) # (!pccount_29))

	.dataa(pccount_29),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[28]~53 ),
	.combout(\pc_count_four_output[29]~54_combout ),
	.cout(\pc_count_four_output[29]~55 ));
// synopsys translate_off
defparam \pc_count_four_output[29]~54 .lut_mask = 16'h5A5F;
defparam \pc_count_four_output[29]~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N22
cycloneive_lcell_comb \branch_count_output[28]~52 (
// Equation(s):
// \branch_count_output[28]~52_combout  = ((temp_npc_28 $ (temp_signZero_16 $ (!\branch_count_output[27]~51 )))) # (GND)
// \branch_count_output[28]~53  = CARRY((temp_npc_28 & ((temp_signZero_16) # (!\branch_count_output[27]~51 ))) # (!temp_npc_28 & (temp_signZero_16 & !\branch_count_output[27]~51 )))

	.dataa(\EXMEM|temp_npc [28]),
	.datab(\EXMEM|temp_signZero [16]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[27]~51 ),
	.combout(\branch_count_output[28]~52_combout ),
	.cout(\branch_count_output[28]~53 ));
// synopsys translate_off
defparam \branch_count_output[28]~52 .lut_mask = 16'h698E;
defparam \branch_count_output[28]~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N24
cycloneive_lcell_comb \branch_count_output[29]~54 (
// Equation(s):
// \branch_count_output[29]~54_combout  = (temp_npc_29 & ((temp_signZero_16 & (\branch_count_output[28]~53  & VCC)) # (!temp_signZero_16 & (!\branch_count_output[28]~53 )))) # (!temp_npc_29 & ((temp_signZero_16 & (!\branch_count_output[28]~53 )) # 
// (!temp_signZero_16 & ((\branch_count_output[28]~53 ) # (GND)))))
// \branch_count_output[29]~55  = CARRY((temp_npc_29 & (!temp_signZero_16 & !\branch_count_output[28]~53 )) # (!temp_npc_29 & ((!\branch_count_output[28]~53 ) # (!temp_signZero_16))))

	.dataa(\EXMEM|temp_npc [29]),
	.datab(\EXMEM|temp_signZero [16]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[28]~53 ),
	.combout(\branch_count_output[29]~54_combout ),
	.cout(\branch_count_output[29]~55 ));
// synopsys translate_off
defparam \branch_count_output[29]~54 .lut_mask = 16'h9617;
defparam \branch_count_output[29]~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N26
cycloneive_lcell_comb \pc_count_four_output[30]~56 (
// Equation(s):
// \pc_count_four_output[30]~56_combout  = (pccount_30 & (\pc_count_four_output[29]~55  $ (GND))) # (!pccount_30 & (!\pc_count_four_output[29]~55  & VCC))
// \pc_count_four_output[30]~57  = CARRY((pccount_30 & !\pc_count_four_output[29]~55 ))

	.dataa(pccount_30),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_count_four_output[29]~55 ),
	.combout(\pc_count_four_output[30]~56_combout ),
	.cout(\pc_count_four_output[30]~57 ));
// synopsys translate_off
defparam \pc_count_four_output[30]~56 .lut_mask = 16'hA50A;
defparam \pc_count_four_output[30]~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N28
cycloneive_lcell_comb \pc_count_four_output[31]~58 (
// Equation(s):
// \pc_count_four_output[31]~58_combout  = \pc_count_four_output[30]~57  $ (pccount_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pccount_31),
	.cin(\pc_count_four_output[30]~57 ),
	.combout(\pc_count_four_output[31]~58_combout ),
	.cout());
// synopsys translate_off
defparam \pc_count_four_output[31]~58 .lut_mask = 16'h0FF0;
defparam \pc_count_four_output[31]~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N26
cycloneive_lcell_comb \branch_count_output[30]~56 (
// Equation(s):
// \branch_count_output[30]~56_combout  = ((temp_npc_30 $ (temp_signZero_16 $ (!\branch_count_output[29]~55 )))) # (GND)
// \branch_count_output[30]~57  = CARRY((temp_npc_30 & ((temp_signZero_16) # (!\branch_count_output[29]~55 ))) # (!temp_npc_30 & (temp_signZero_16 & !\branch_count_output[29]~55 )))

	.dataa(\EXMEM|temp_npc [30]),
	.datab(\EXMEM|temp_signZero [16]),
	.datac(gnd),
	.datad(vcc),
	.cin(\branch_count_output[29]~55 ),
	.combout(\branch_count_output[30]~56_combout ),
	.cout(\branch_count_output[30]~57 ));
// synopsys translate_off
defparam \branch_count_output[30]~56 .lut_mask = 16'h698E;
defparam \branch_count_output[30]~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N28
cycloneive_lcell_comb \branch_count_output[31]~58 (
// Equation(s):
// \branch_count_output[31]~58_combout  = temp_npc_31 $ (\branch_count_output[30]~57  $ (temp_signZero_16))

	.dataa(\EXMEM|temp_npc [31]),
	.datab(gnd),
	.datac(gnd),
	.datad(\EXMEM|temp_signZero [16]),
	.cin(\branch_count_output[30]~57 ),
	.combout(\branch_count_output[31]~58_combout ),
	.cout());
// synopsys translate_off
defparam \branch_count_output[31]~58 .lut_mask = 16'hA55A;
defparam \branch_count_output[31]~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: DDIOOUTCELL_X58_Y73_N25
dffeas \dpif.halt (
	.clk(CPUCLK),
	.d(\EXMEM|temp_halt_out~q ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dpifhalt),
	.prn(vcc));
// synopsys translate_off
defparam \dpif.halt .is_wysiwyg = "true";
defparam \dpif.halt .power_up = "low";
// synopsys translate_on

endmodule

module alu (
	temp_ALUop_output_0,
	temp_imemload_output_7,
	temp_ALUsrc_output_1,
	temp_ALUsrc_output_0,
	Mux30,
	alu_b_mux_output_1,
	alu_b_mux_output_11,
	Mux16,
	Mux301,
	alu_a_mux_output_1,
	temp_ALUop_output_1,
	alu_b_mux_output_0,
	temp_imemload_output_6,
	Mux31,
	alu_b_mux_output_01,
	alu_a_mux_output_0,
	alu_a_mux_output_2,
	Mux311,
	alu_a_mux_output_4,
	alu_a_mux_output_3,
	alu_a_mux_output_31,
	Mux29,
	alu_b_mux_output_2,
	Mux291,
	alu_a_mux_output_8,
	alu_a_mux_output_7,
	alu_a_mux_output_6,
	alu_a_mux_output_5,
	Mux28,
	alu_b_mux_output_3,
	Mux281,
	alu_a_mux_output_16,
	alu_a_mux_output_14,
	alu_a_mux_output_15,
	alu_a_mux_output_13,
	alu_a_mux_output_12,
	alu_a_mux_output_10,
	alu_a_mux_output_11,
	alu_a_mux_output_9,
	Mux27,
	alu_b_mux_output_4,
	Mux271,
	alu_a_mux_output_311,
	alu_a_mux_output_30,
	alu_a_mux_output_29,
	alu_a_mux_output_26,
	alu_a_mux_output_25,
	alu_a_mux_output_28,
	alu_a_mux_output_27,
	alu_a_mux_output_17,
	alu_a_mux_output_20,
	alu_a_mux_output_19,
	alu_a_mux_output_18,
	alu_a_mux_output_24,
	alu_a_mux_output_23,
	alu_a_mux_output_22,
	alu_a_mux_output_21,
	Mux161,
	Mux19,
	Mux4,
	Mux13,
	Mux14,
	Mux15,
	Mux0,
	Mux1,
	Mux2,
	Mux3,
	Mux5,
	Mux6,
	Mux7,
	Mux8,
	Mux9,
	Mux10,
	Mux11,
	Mux12,
	Mux17,
	Mux21,
	alu_b_mux_output_14,
	Mux22,
	Mux23,
	alu_b_mux_output_7,
	Mux24,
	alu_b_mux_output_6,
	Mux25,
	alu_b_mux_output_5,
	temp_imemload_output_5,
	Mux26,
	Mux18,
	Mux20,
	temp_ALUop_output_2,
	temp_ALUop_output_3,
	Mux302,
	Mux171,
	Mux312,
	Mux292,
	Mux282,
	alu_a_mux_output_32,
	Mux261,
	Mux272,
	Mux241,
	Mux251,
	Mux221,
	Mux222,
	Mux191,
	Mux231,
	Mux232,
	Mux201,
	Mux202,
	Mux211,
	Mux212,
	Mux181,
	Mux182,
	Mux192,
	Mux193,
	Mux162,
	Mux163,
	Mux172,
	Mux173,
	Mux141,
	Mux142,
	Mux151,
	Mux152,
	Mux121,
	Mux122,
	Mux131,
	Mux132,
	Mux111,
	Mux112,
	Mux101,
	Mux102,
	Mux81,
	Mux82,
	Mux91,
	Mux92,
	Mux61,
	Mux41,
	Mux210,
	Mux32,
	Mux01,
	Mux02,
	Mux110,
	Equal0,
	Mux113,
	Mux51,
	Mux71,
	devpor,
	devclrn,
	devoe);
input 	temp_ALUop_output_0;
input 	temp_imemload_output_7;
input 	temp_ALUsrc_output_1;
input 	temp_ALUsrc_output_0;
input 	Mux30;
input 	alu_b_mux_output_1;
input 	alu_b_mux_output_11;
input 	Mux16;
input 	Mux301;
input 	alu_a_mux_output_1;
input 	temp_ALUop_output_1;
input 	alu_b_mux_output_0;
input 	temp_imemload_output_6;
input 	Mux31;
input 	alu_b_mux_output_01;
input 	alu_a_mux_output_0;
input 	alu_a_mux_output_2;
input 	Mux311;
input 	alu_a_mux_output_4;
input 	alu_a_mux_output_3;
input 	alu_a_mux_output_31;
input 	Mux29;
input 	alu_b_mux_output_2;
input 	Mux291;
input 	alu_a_mux_output_8;
input 	alu_a_mux_output_7;
input 	alu_a_mux_output_6;
input 	alu_a_mux_output_5;
input 	Mux28;
input 	alu_b_mux_output_3;
input 	Mux281;
input 	alu_a_mux_output_16;
input 	alu_a_mux_output_14;
input 	alu_a_mux_output_15;
input 	alu_a_mux_output_13;
input 	alu_a_mux_output_12;
input 	alu_a_mux_output_10;
input 	alu_a_mux_output_11;
input 	alu_a_mux_output_9;
input 	Mux27;
input 	alu_b_mux_output_4;
input 	Mux271;
input 	alu_a_mux_output_311;
input 	alu_a_mux_output_30;
input 	alu_a_mux_output_29;
input 	alu_a_mux_output_26;
input 	alu_a_mux_output_25;
input 	alu_a_mux_output_28;
input 	alu_a_mux_output_27;
input 	alu_a_mux_output_17;
input 	alu_a_mux_output_20;
input 	alu_a_mux_output_19;
input 	alu_a_mux_output_18;
input 	alu_a_mux_output_24;
input 	alu_a_mux_output_23;
input 	alu_a_mux_output_22;
input 	alu_a_mux_output_21;
input 	Mux161;
input 	Mux19;
input 	Mux4;
input 	Mux13;
input 	Mux14;
input 	Mux15;
input 	Mux0;
input 	Mux1;
input 	Mux2;
input 	Mux3;
input 	Mux5;
input 	Mux6;
input 	Mux7;
input 	Mux8;
input 	Mux9;
input 	Mux10;
input 	Mux11;
input 	Mux12;
input 	Mux17;
input 	Mux21;
input 	alu_b_mux_output_14;
input 	Mux22;
input 	Mux23;
input 	alu_b_mux_output_7;
input 	Mux24;
input 	alu_b_mux_output_6;
input 	Mux25;
input 	alu_b_mux_output_5;
input 	temp_imemload_output_5;
input 	Mux26;
input 	Mux18;
input 	Mux20;
input 	temp_ALUop_output_2;
input 	temp_ALUop_output_3;
output 	Mux302;
input 	Mux171;
output 	Mux312;
output 	Mux292;
output 	Mux282;
input 	alu_a_mux_output_32;
output 	Mux261;
output 	Mux272;
output 	Mux241;
output 	Mux251;
output 	Mux221;
output 	Mux222;
output 	Mux191;
output 	Mux231;
output 	Mux232;
output 	Mux201;
output 	Mux202;
output 	Mux211;
output 	Mux212;
output 	Mux181;
output 	Mux182;
output 	Mux192;
output 	Mux193;
output 	Mux162;
output 	Mux163;
output 	Mux172;
output 	Mux173;
output 	Mux141;
output 	Mux142;
output 	Mux151;
output 	Mux152;
output 	Mux121;
output 	Mux122;
output 	Mux131;
output 	Mux132;
output 	Mux111;
output 	Mux112;
output 	Mux101;
output 	Mux102;
output 	Mux81;
output 	Mux82;
output 	Mux91;
output 	Mux92;
output 	Mux61;
output 	Mux41;
output 	Mux210;
output 	Mux32;
output 	Mux01;
output 	Mux02;
output 	Mux110;
output 	Equal0;
output 	Mux113;
output 	Mux51;
output 	Mux71;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add0~8_combout ;
wire \Add0~13_combout ;
wire \Add0~16_combout ;
wire \Add0~4_combout ;
wire \ShiftRight0~2_combout ;
wire \ShiftRight0~3_combout ;
wire \ShiftRight0~4_combout ;
wire \ShiftRight0~5_combout ;
wire \ShiftRight0~7_combout ;
wire \ShiftRight0~8_combout ;
wire \ShiftRight0~16_combout ;
wire \ShiftLeft0~5_combout ;
wire \ShiftRight0~29_combout ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux31~3_combout ;
wire \ShiftRight0~30_combout ;
wire \ShiftRight0~32_combout ;
wire \ShiftRight0~36_combout ;
wire \ShiftRight0~42_combout ;
wire \ShiftRight0~50_combout ;
wire \ShiftRight0~52_combout ;
wire \Mux31~4_combout ;
wire \Mux31~5_combout ;
wire \ShiftRight0~63_combout ;
wire \ShiftRight0~69_combout ;
wire \ShiftRight0~70_combout ;
wire \ShiftLeft0~19_combout ;
wire \OUTPUT~0_combout ;
wire \Mux29~6_combout ;
wire \OUTPUT~1_combout ;
wire \Mux26~2_combout ;
wire \ShiftLeft0~27_combout ;
wire \Mux24~0_combout ;
wire \ShiftLeft0~38_combout ;
wire \ShiftLeft0~42_combout ;
wire \Mux20~1_combout ;
wire \ShiftRight0~106_combout ;
wire \Mux19~8_combout ;
wire \ShiftLeft0~75_combout ;
wire \Mux12~4_combout ;
wire \Mux13~1_combout ;
wire \Mux7~0_combout ;
wire \ShiftLeft0~99_combout ;
wire \ShiftLeft0~100_combout ;
wire \ShiftLeft0~101_combout ;
wire \Mux4~2_combout ;
wire \ShiftLeft0~103_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \OUTPUT~3_combout ;
wire \Mux10~6_combout ;
wire \Equal0~15_combout ;
wire \Equal0~16_combout ;
wire \Equal0~18_combout ;
wire \Add0~105_combout ;
wire \Mux2~15_combout ;
wire \ShiftLeft0~13_combout ;
wire \ShiftLeft0~12_combout ;
wire \ShiftLeft0~14_combout ;
wire \ShiftLeft0~15_combout ;
wire \Mux30~2_combout ;
wire \Mux30~3_combout ;
wire \Add0~106_combout ;
wire \Add0~5_combout ;
wire \Add0~7_cout ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~17_cout ;
wire \LessThan0~19_cout ;
wire \LessThan0~21_cout ;
wire \LessThan0~23_cout ;
wire \LessThan0~25_cout ;
wire \LessThan0~27_cout ;
wire \LessThan0~29_cout ;
wire \LessThan0~31_cout ;
wire \LessThan0~33_cout ;
wire \LessThan0~35_cout ;
wire \LessThan0~37_cout ;
wire \LessThan0~39_cout ;
wire \LessThan0~41_cout ;
wire \LessThan0~43_cout ;
wire \LessThan0~45_cout ;
wire \LessThan0~47_cout ;
wire \LessThan0~49_cout ;
wire \LessThan0~51_cout ;
wire \LessThan0~53_cout ;
wire \LessThan0~55_cout ;
wire \LessThan0~57_cout ;
wire \LessThan0~59_cout ;
wire \LessThan0~61_cout ;
wire \LessThan0~62_combout ;
wire \LessThan1~1_cout ;
wire \LessThan1~3_cout ;
wire \LessThan1~5_cout ;
wire \LessThan1~7_cout ;
wire \LessThan1~9_cout ;
wire \LessThan1~11_cout ;
wire \LessThan1~13_cout ;
wire \LessThan1~15_cout ;
wire \LessThan1~17_cout ;
wire \LessThan1~19_cout ;
wire \LessThan1~21_cout ;
wire \LessThan1~23_cout ;
wire \LessThan1~25_cout ;
wire \LessThan1~27_cout ;
wire \LessThan1~29_cout ;
wire \LessThan1~31_cout ;
wire \LessThan1~33_cout ;
wire \LessThan1~35_cout ;
wire \LessThan1~37_cout ;
wire \LessThan1~39_cout ;
wire \LessThan1~41_cout ;
wire \LessThan1~43_cout ;
wire \LessThan1~45_cout ;
wire \LessThan1~47_cout ;
wire \LessThan1~49_cout ;
wire \LessThan1~51_cout ;
wire \LessThan1~53_cout ;
wire \LessThan1~55_cout ;
wire \LessThan1~57_cout ;
wire \LessThan1~59_cout ;
wire \LessThan1~61_cout ;
wire \LessThan1~62_combout ;
wire \Mux31~2_combout ;
wire \Mux31~6_combout ;
wire \Mux31~7_combout ;
wire \Mux31~8_combout ;
wire \Mux29~11_combout ;
wire \Mux19~1_combout ;
wire \Mux29~0_combout ;
wire \ShiftRight0~34_combout ;
wire \ShiftRight0~57_combout ;
wire \ShiftRight0~56_combout ;
wire \ShiftRight0~58_combout ;
wire \ShiftRight0~31_combout ;
wire \Mux29~1_combout ;
wire \Mux29~2_combout ;
wire \ShiftRight0~71_combout ;
wire \ShiftRight0~72_combout ;
wire \ShiftRight0~73_combout ;
wire \ShiftRight0~65_combout ;
wire \ShiftRight0~66_combout ;
wire \ShiftRight0~67_combout ;
wire \ShiftRight0~44_combout ;
wire \ShiftRight0~68_combout ;
wire \ShiftRight0~74_combout ;
wire \Mux29~3_combout ;
wire \Mux29~7_combout ;
wire \Mux19~2_combout ;
wire \ShiftLeft0~9_combout ;
wire \ShiftLeft0~10_combout ;
wire \ShiftLeft0~4_combout ;
wire \ShiftLeft0~2_combout ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~6_combout ;
wire \ShiftLeft0~7_combout ;
wire \ShiftLeft0~11_combout ;
wire \Mux29~8_combout ;
wire \Mux29~9_combout ;
wire \Mux29~10_combout ;
wire \ShiftRight0~37_combout ;
wire \ShiftRight0~60_combout ;
wire \ShiftRight0~76_combout ;
wire \ShiftRight0~77_combout ;
wire \ShiftRight0~78_combout ;
wire \ShiftRight0~79_combout ;
wire \ShiftRight0~6_combout ;
wire \ShiftRight0~59_combout ;
wire \ShiftRight0~39_combout ;
wire \ShiftRight0~75_combout ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \Mux29~5_combout ;
wire \ShiftLeft0~20_combout ;
wire \ShiftLeft0~21_combout ;
wire \ShiftLeft0~8_combout ;
wire \Mux19~0_combout ;
wire \Mux29~4_combout ;
wire \Mux28~2_combout ;
wire \Mux28~3_combout ;
wire \Mux28~4_combout ;
wire \Mux28~5_combout ;
wire \Mux26~5_combout ;
wire \Add0~18_combout ;
wire \Add0~19_combout ;
wire \Add0~20_combout ;
wire \Add0~15_combout ;
wire \Add0~12_combout ;
wire \Add0~11 ;
wire \Add0~14 ;
wire \Add0~17 ;
wire \Add0~22 ;
wire \Add0~23_combout ;
wire \Mux27~3_combout ;
wire \Mux27~2_combout ;
wire \ShiftRight0~23_combout ;
wire \Mux1~0_combout ;
wire \ShiftRight0~24_combout ;
wire \ShiftRight0~10_combout ;
wire \ShiftRight0~9_combout ;
wire \ShiftRight0~11_combout ;
wire \ShiftRight0~90_combout ;
wire \Mux26~0_combout ;
wire \ShiftRight0~19_combout ;
wire \ShiftRight0~20_combout ;
wire \ShiftRight0~26_combout ;
wire \ShiftRight0~91_combout ;
wire \ShiftRight0~92_combout ;
wire \ShiftRight0~12_combout ;
wire \ShiftRight0~13_combout ;
wire \ShiftRight0~14_combout ;
wire \Mux26~1_combout ;
wire \ShiftLeft0~26_combout ;
wire \Mux27~4_combout ;
wire \Mux26~3_combout ;
wire \Mux26~4_combout ;
wire \Mux27~12_combout ;
wire \Mux27~10_combout ;
wire \Add0~21_combout ;
wire \ShiftRight0~53_combout ;
wire \ShiftRight0~54_combout ;
wire \ShiftRight0~46_combout ;
wire \ShiftRight0~94_combout ;
wire \ShiftRight0~43_combout ;
wire \ShiftRight0~45_combout ;
wire \ShiftRight0~95_combout ;
wire \ShiftRight0~40_combout ;
wire \ShiftRight0~33_combout ;
wire \ShiftRight0~35_combout ;
wire \Mux27~5_combout ;
wire \Mux27~6_combout ;
wire \ShiftLeft0~22_combout ;
wire \ShiftLeft0~28_combout ;
wire \ShiftLeft0~16_combout ;
wire \ShiftLeft0~29_combout ;
wire \Mux27~7_combout ;
wire \Mux27~8_combout ;
wire \Mux27~9_combout ;
wire \Mux24~5_combout ;
wire \ShiftRight0~80_combout ;
wire \ShiftRight0~82_combout ;
wire \ShiftRight0~81_combout ;
wire \ShiftRight0~97_combout ;
wire \ShiftRight0~98_combout ;
wire \Mux24~1_combout ;
wire \ShiftLeft0~32_combout ;
wire \ShiftLeft0~31_combout ;
wire \ShiftLeft0~33_combout ;
wire \ShiftLeft0~30_combout ;
wire \ShiftLeft0~34_combout ;
wire \Mux24~2_combout ;
wire \Mux24~3_combout ;
wire \Mux24~4_combout ;
wire \Add0~25_combout ;
wire \Add0~26_combout ;
wire \Add0~27_combout ;
wire \Add0~28_combout ;
wire \Add0~24 ;
wire \Add0~30 ;
wire \Add0~31_combout ;
wire \Add0~29_combout ;
wire \Mux25~5_combout ;
wire \ShiftLeft0~18_combout ;
wire \ShiftLeft0~104_combout ;
wire \ShiftLeft0~23_combout ;
wire \ShiftLeft0~35_combout ;
wire \ShiftLeft0~36_combout ;
wire \Mux25~2_combout ;
wire \ShiftRight0~61_combout ;
wire \Mux25~0_combout ;
wire \ShiftRight0~99_combout ;
wire \ShiftRight0~62_combout ;
wire \ShiftRight0~100_combout ;
wire \ShiftRight0~101_combout ;
wire \ShiftRight0~102_combout ;
wire \Mux25~1_combout ;
wire \Mux25~3_combout ;
wire \Mux25~4_combout ;
wire \ShiftRight0~15_combout ;
wire \Mux19~3_combout ;
wire \ShiftRight0~25_combout ;
wire \ShiftRight0~27_combout ;
wire \ShiftLeft0~37_combout ;
wire \ShiftLeft0~39_combout ;
wire \ShiftLeft0~24_combout ;
wire \ShiftLeft0~40_combout ;
wire \ShiftLeft0~41_combout ;
wire \Mux22~1_combout ;
wire \Mux19~4_combout ;
wire \Mux19~5_combout ;
wire \Mux22~2_combout ;
wire \Mux22~3_combout ;
wire \Add0~33_combout ;
wire \Add0~34_combout ;
wire \Add0~32 ;
wire \Add0~36 ;
wire \Add0~37_combout ;
wire \Mux22~4_combout ;
wire \Add0~35_combout ;
wire \Mux23~4_combout ;
wire \ShiftRight0~38_combout ;
wire \ShiftRight0~41_combout ;
wire \ShiftRight0~47_combout ;
wire \ShiftRight0~48_combout ;
wire \ShiftRight0~49_combout ;
wire \ShiftRight0~51_combout ;
wire \ShiftLeft0~43_combout ;
wire \ShiftLeft0~44_combout ;
wire \ShiftLeft0~45_combout ;
wire \Mux23~1_combout ;
wire \Mux23~2_combout ;
wire \Mux23~3_combout ;
wire \Mux20~4_combout ;
wire \Add0~39_combout ;
wire \Add0~40_combout ;
wire \Add0~38 ;
wire \Add0~42 ;
wire \Add0~43_combout ;
wire \ShiftRight0~83_combout ;
wire \ShiftRight0~105_combout ;
wire \Mux20~2_combout ;
wire \ShiftRight0~84_combout ;
wire \ShiftRight0~85_combout ;
wire \ShiftRight0~86_combout ;
wire \ShiftRight0~87_combout ;
wire \ShiftRight0~88_combout ;
wire \Mux20~3_combout ;
wire \ShiftRight0~64_combout ;
wire \ShiftLeft0~46_combout ;
wire \ShiftLeft0~51_combout ;
wire \ShiftLeft0~52_combout ;
wire \ShiftLeft0~53_combout ;
wire \Mux21~1_combout ;
wire \Mux21~2_combout ;
wire \Mux21~3_combout ;
wire \Mux21~4_combout ;
wire \Add0~41_combout ;
wire \Add0~45_combout ;
wire \Add0~44 ;
wire \Add0~48 ;
wire \Add0~49_combout ;
wire \ShiftLeft0~55_combout ;
wire \ShiftLeft0~54_combout ;
wire \ShiftLeft0~56_combout ;
wire \ShiftLeft0~57_combout ;
wire \ShiftLeft0~25_combout ;
wire \ShiftLeft0~58_combout ;
wire \Mux18~1_combout ;
wire \ShiftRight0~17_combout ;
wire \ShiftRight0~18_combout ;
wire \ShiftRight0~111_combout ;
wire \Mux18~2_combout ;
wire \Mux18~3_combout ;
wire \Mux18~4_combout ;
wire \Add0~46_combout ;
wire \Add0~47_combout ;
wire \Mux19~11_combout ;
wire \ShiftRight0~93_combout ;
wire \ShiftRight0~108_combout ;
wire \Mux19~9_combout ;
wire \Mux19~10_combout ;
wire \Mux16~4_combout ;
wire \Add0~51_combout ;
wire \Add0~50 ;
wire \Add0~54 ;
wire \Add0~55_combout ;
wire \ShiftLeft0~47_combout ;
wire \ShiftLeft0~48_combout ;
wire \ShiftLeft0~65_combout ;
wire \Mux16~1_combout ;
wire \Mux16~2_combout ;
wire \ShiftRight0~96_combout ;
wire \Mux16~3_combout ;
wire \Add0~52_combout ;
wire \Add0~53_combout ;
wire \Mux17~4_combout ;
wire \ShiftRight0~110_combout ;
wire \ShiftLeft0~62_combout ;
wire \ShiftLeft0~66_combout ;
wire \ShiftLeft0~67_combout ;
wire \Mux17~1_combout ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \ShiftLeft0~70_combout ;
wire \Mux12~2_combout ;
wire \ShiftRight0~21_combout ;
wire \ShiftRight0~28_combout ;
wire \Mux14~1_combout ;
wire \Mux12~0_combout ;
wire \Mux14~2_combout ;
wire \Mux14~3_combout ;
wire \Add0~57_combout ;
wire \Add0~56 ;
wire \Add0~60 ;
wire \Add0~61_combout ;
wire \Add0~58_combout ;
wire \Add0~59_combout ;
wire \ShiftRight0~55_combout ;
wire \ShiftLeft0~17_combout ;
wire \Mux15~1_combout ;
wire \ShiftLeft0~59_combout ;
wire \ShiftLeft0~72_combout ;
wire \ShiftLeft0~73_combout ;
wire \Mux15~2_combout ;
wire \Mux15~3_combout ;
wire \Add0~63_combout ;
wire \Add0~62 ;
wire \Add0~66 ;
wire \Add0~67_combout ;
wire \ShiftLeft0~49_combout ;
wire \ShiftLeft0~74_combout ;
wire \ShiftLeft0~63_combout ;
wire \ShiftLeft0~64_combout ;
wire \ShiftLeft0~76_combout ;
wire \ShiftRight0~89_combout ;
wire \Mux12~1_combout ;
wire \Mux12~5_combout ;
wire \Mux12~6_combout ;
wire \Mux12~7_combout ;
wire \Mux13~4_combout ;
wire \ShiftLeft0~78_combout ;
wire \ShiftLeft0~77_combout ;
wire \ShiftLeft0~79_combout ;
wire \Mux13~2_combout ;
wire \Mux13~3_combout ;
wire \Add0~64_combout ;
wire \Add0~65_combout ;
wire \ShiftLeft0~60_combout ;
wire \ShiftLeft0~80_combout ;
wire \ShiftLeft0~81_combout ;
wire \ShiftLeft0~71_combout ;
wire \ShiftLeft0~82_combout ;
wire \Mux11~1_combout ;
wire \Mux11~2_combout ;
wire \Mux11~3_combout ;
wire \Add0~69_combout ;
wire \Add0~68 ;
wire \Add0~70_combout ;
wire \Mux11~4_combout ;
wire \Add0~72_combout ;
wire \Add0~71 ;
wire \Add0~73_combout ;
wire \ShiftLeft0~83_combout ;
wire \ShiftLeft0~84_combout ;
wire \ShiftLeft0~68_combout ;
wire \ShiftRight0~22_combout ;
wire \ShiftLeft0~69_combout ;
wire \ShiftLeft0~85_combout ;
wire \Mux10~1_combout ;
wire \Mux10~2_combout ;
wire \Mux10~3_combout ;
wire \Mux10~4_combout ;
wire \Mux8~4_combout ;
wire \ShiftLeft0~86_combout ;
wire \ShiftLeft0~87_combout ;
wire \ShiftLeft0~88_combout ;
wire \Mux8~1_combout ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \Add0~75_combout ;
wire \Add0~76_combout ;
wire \Add0~74 ;
wire \Add0~78 ;
wire \Add0~79_combout ;
wire \Mux9~4_combout ;
wire \ShiftLeft0~89_combout ;
wire \ShiftLeft0~90_combout ;
wire \ShiftLeft0~91_combout ;
wire \Mux9~1_combout ;
wire \Mux9~2_combout ;
wire \Mux9~3_combout ;
wire \Add0~77_combout ;
wire \Mux6~6_combout ;
wire \ShiftLeft0~92_combout ;
wire \ShiftLeft0~93_combout ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \Mux6~8_combout ;
wire \ShiftRight0~103_combout ;
wire \Mux6~4_combout ;
wire \Mux6~5_combout ;
wire \Add0~81_combout ;
wire \Add0~82_combout ;
wire \Add0~80 ;
wire \Add0~84 ;
wire \Add0~85_combout ;
wire \ShiftLeft0~50_combout ;
wire \Mux4~3_combout ;
wire \Mux4~8_combout ;
wire \Mux4~4_combout ;
wire \Mux4~5_combout ;
wire \Add0~90_combout ;
wire \Add0~86 ;
wire \Add0~89 ;
wire \Add0~91_combout ;
wire \Mux4~6_combout ;
wire \ShiftLeft0~102_combout ;
wire \Mux2~3_combout ;
wire \Mux2~4_combout ;
wire \Mux2~6_combout ;
wire \OUTPUT~2_combout ;
wire \Mux2~7_combout ;
wire \Mux2~8_combout ;
wire \Mux2~9_combout ;
wire \Mux2~10_combout ;
wire \Mux2~11_combout ;
wire \Mux2~12_combout ;
wire \Mux2~13_combout ;
wire \Add0~93_combout ;
wire \Add0~92 ;
wire \Add0~96 ;
wire \Add0~97_combout ;
wire \Mux2~5_combout ;
wire \Mux3~2_combout ;
wire \Mux2~2_combout ;
wire \ShiftLeft0~61_combout ;
wire \Mux3~3_combout ;
wire \Mux3~4_combout ;
wire \Mux3~5_combout ;
wire \Mux3~6_combout ;
wire \Mux3~7_combout ;
wire \Mux3~8_combout ;
wire \Add0~94_combout ;
wire \Add0~95_combout ;
wire \Add0~99_combout ;
wire \Add0~98 ;
wire \Add0~102 ;
wire \Add0~103_combout ;
wire \ShiftRight0~109_combout ;
wire \Mux0~3_combout ;
wire \Mux0~4_combout ;
wire \Mux1~1_combout ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux0~5_combout ;
wire \Mux0~6_combout ;
wire \Equal0~4_combout ;
wire \Equal0~5_combout ;
wire \Mux9~6_combout ;
wire \Mux11~6_combout ;
wire \Equal0~2_combout ;
wire \Equal0~3_combout ;
wire \Equal0~6_combout ;
wire \Equal0~7_combout ;
wire \Equal0~8_combout ;
wire \Equal0~9_combout ;
wire \Mux1~8_combout ;
wire \Equal0~10_combout ;
wire \Mux23~6_combout ;
wire \Mux22~6_combout ;
wire \Mux14~5_combout ;
wire \Mux16~6_combout ;
wire \Mux18~6_combout ;
wire \Equal0~11_combout ;
wire \Equal0~12_combout ;
wire \Equal0~13_combout ;
wire \Mux13~6_combout ;
wire \Mux8~6_combout ;
wire \Mux12~9_combout ;
wire \Equal0~14_combout ;
wire \Equal0~17_combout ;
wire \Equal0~19_combout ;
wire \Equal0~23_combout ;
wire \Equal0~20_combout ;
wire \Equal0~21_combout ;
wire \Mux1~3_combout ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux1~6_combout ;
wire \Mux1~7_combout ;
wire \Mux1~9_combout ;
wire \Add0~100_combout ;
wire \Add0~101_combout ;
wire \Mux5~7_combout ;
wire \ShiftRight0~107_combout ;
wire \ShiftLeft0~96_combout ;
wire \ShiftLeft0~97_combout ;
wire \ShiftLeft0~98_combout ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \Mux5~6_combout ;
wire \Mux5~4_combout ;
wire \Mux5~5_combout ;
wire \Add0~87_combout ;
wire \Add0~88_combout ;
wire \ShiftRight0~104_combout ;
wire \ShiftLeft0~94_combout ;
wire \ShiftLeft0~95_combout ;
wire \Mux7~1_combout ;
wire \Mux7~2_combout ;
wire \Mux7~3_combout ;
wire \Mux7~4_combout ;
wire \Mux7~5_combout ;
wire \Mux7~6_combout ;
wire \Add0~83_combout ;


// Location: LCCOMB_X67_Y42_N18
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = (alu_a_mux_output_0 & ((\Add0~5_combout  & (\Add0~7_cout  & VCC)) # (!\Add0~5_combout  & (!\Add0~7_cout )))) # (!alu_a_mux_output_0 & ((\Add0~5_combout  & (!\Add0~7_cout )) # (!\Add0~5_combout  & ((\Add0~7_cout ) # (GND)))))
// \Add0~9  = CARRY((alu_a_mux_output_0 & (!\Add0~5_combout  & !\Add0~7_cout )) # (!alu_a_mux_output_0 & ((!\Add0~7_cout ) # (!\Add0~5_combout ))))

	.dataa(alu_a_mux_output_0),
	.datab(\Add0~5_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7_cout ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'h9617;
defparam \Add0~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N22
cycloneive_lcell_comb \Add0~13 (
// Equation(s):
// \Add0~13_combout  = (alu_a_mux_output_2 & ((\Add0~12_combout  & (\Add0~11  & VCC)) # (!\Add0~12_combout  & (!\Add0~11 )))) # (!alu_a_mux_output_2 & ((\Add0~12_combout  & (!\Add0~11 )) # (!\Add0~12_combout  & ((\Add0~11 ) # (GND)))))
// \Add0~14  = CARRY((alu_a_mux_output_2 & (!\Add0~12_combout  & !\Add0~11 )) # (!alu_a_mux_output_2 & ((!\Add0~11 ) # (!\Add0~12_combout ))))

	.dataa(alu_a_mux_output_2),
	.datab(\Add0~12_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~13_combout ),
	.cout(\Add0~14 ));
// synopsys translate_off
defparam \Add0~13 .lut_mask = 16'h9617;
defparam \Add0~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N24
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = ((alu_a_mux_output_31 $ (\Add0~15_combout  $ (!\Add0~14 )))) # (GND)
// \Add0~17  = CARRY((alu_a_mux_output_31 & ((\Add0~15_combout ) # (!\Add0~14 ))) # (!alu_a_mux_output_31 & (\Add0~15_combout  & !\Add0~14 )))

	.dataa(alu_a_mux_output_31),
	.datab(\Add0~15_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~14 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'h698E;
defparam \Add0~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N4
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = temp_ALUop_output_0 $ ((((!Mux16 & alu_b_mux_output_11)) # (!\Add0~105_combout )))

	.dataa(Mux16),
	.datab(\Add0~105_combout ),
	.datac(temp_ALUop_output_0),
	.datad(alu_b_mux_output_11),
	.cin(gnd),
	.combout(\Add0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'h87C3;
defparam \Add0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N4
cycloneive_lcell_comb \ShiftRight0~2 (
// Equation(s):
// \ShiftRight0~2_combout  = (!Mux301 & ((Mux311 & ((alu_a_mux_output_2))) # (!Mux311 & (alu_a_mux_output_1))))

	.dataa(Mux301),
	.datab(Mux311),
	.datac(alu_a_mux_output_1),
	.datad(alu_a_mux_output_2),
	.cin(gnd),
	.combout(\ShiftRight0~2_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~2 .lut_mask = 16'h5410;
defparam \ShiftRight0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N10
cycloneive_lcell_comb \ShiftRight0~3 (
// Equation(s):
// \ShiftRight0~3_combout  = (Mux311 & ((alu_a_mux_output_4))) # (!Mux311 & (alu_a_mux_output_31))

	.dataa(alu_a_mux_output_31),
	.datab(gnd),
	.datac(alu_a_mux_output_4),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftRight0~3_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~3 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N8
cycloneive_lcell_comb \ShiftRight0~4 (
// Equation(s):
// \ShiftRight0~4_combout  = (!Mux291 & ((\ShiftRight0~2_combout ) # ((\ShiftRight0~3_combout  & Mux301))))

	.dataa(\ShiftRight0~3_combout ),
	.datab(Mux291),
	.datac(\ShiftRight0~2_combout ),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftRight0~4_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~4 .lut_mask = 16'h3230;
defparam \ShiftRight0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N24
cycloneive_lcell_comb \ShiftRight0~5 (
// Equation(s):
// \ShiftRight0~5_combout  = (Mux301 & ((Mux311 & ((alu_a_mux_output_8))) # (!Mux311 & (alu_a_mux_output_7))))

	.dataa(Mux311),
	.datab(Mux301),
	.datac(alu_a_mux_output_7),
	.datad(alu_a_mux_output_8),
	.cin(gnd),
	.combout(\ShiftRight0~5_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~5 .lut_mask = 16'hC840;
defparam \ShiftRight0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N12
cycloneive_lcell_comb \ShiftRight0~7 (
// Equation(s):
// \ShiftRight0~7_combout  = (\ShiftRight0~5_combout ) # ((!Mux301 & \ShiftRight0~6_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~5_combout ),
	.datac(Mux301),
	.datad(\ShiftRight0~6_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~7 .lut_mask = 16'hCFCC;
defparam \ShiftRight0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N20
cycloneive_lcell_comb \ShiftRight0~8 (
// Equation(s):
// \ShiftRight0~8_combout  = (!Mux281 & ((\ShiftRight0~4_combout ) # ((\ShiftRight0~7_combout  & Mux291))))

	.dataa(\ShiftRight0~7_combout ),
	.datab(Mux281),
	.datac(Mux291),
	.datad(\ShiftRight0~4_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~8 .lut_mask = 16'h3320;
defparam \ShiftRight0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N22
cycloneive_lcell_comb \ShiftRight0~16 (
// Equation(s):
// \ShiftRight0~16_combout  = (!Mux271 & ((\ShiftRight0~8_combout ) # ((\ShiftRight0~15_combout  & Mux281))))

	.dataa(\ShiftRight0~15_combout ),
	.datab(\ShiftRight0~8_combout ),
	.datac(Mux271),
	.datad(Mux281),
	.cin(gnd),
	.combout(\ShiftRight0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~16 .lut_mask = 16'h0E0C;
defparam \ShiftRight0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N30
cycloneive_lcell_comb \ShiftLeft0~5 (
// Equation(s):
// \ShiftLeft0~5_combout  = (Mux9) # ((Mux10) # ((Mux11) # (Mux12)))

	.dataa(Mux9),
	.datab(Mux10),
	.datac(Mux11),
	.datad(Mux12),
	.cin(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~5 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N30
cycloneive_lcell_comb \ShiftRight0~29 (
// Equation(s):
// \ShiftRight0~29_combout  = (!\ShiftLeft0~11_combout  & ((\ShiftRight0~16_combout ) # ((Mux271 & \ShiftRight0~28_combout ))))

	.dataa(Mux271),
	.datab(\ShiftRight0~28_combout ),
	.datac(\ShiftRight0~16_combout ),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~29 .lut_mask = 16'h00F8;
defparam \ShiftRight0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N22
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (!temp_ALUop_output_1 & ((Mux311 & (!alu_a_mux_output_0 & !temp_ALUop_output_0)) # (!Mux311 & (alu_a_mux_output_0 $ (temp_ALUop_output_0)))))

	.dataa(Mux311),
	.datab(alu_a_mux_output_0),
	.datac(temp_ALUop_output_0),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'h0016;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N12
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (\Mux31~0_combout ) # ((temp_ALUop_output_1 & \Add0~8_combout ))

	.dataa(gnd),
	.datab(temp_ALUop_output_1),
	.datac(\Mux31~0_combout ),
	.datad(\Add0~8_combout ),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hFCF0;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N6
cycloneive_lcell_comb \Mux31~3 (
// Equation(s):
// \Mux31~3_combout  = (temp_ALUop_output_1 & (((alu_a_mux_output_0) # (Mux311)))) # (!temp_ALUop_output_1 & (Mux271))

	.dataa(Mux271),
	.datab(alu_a_mux_output_0),
	.datac(Mux311),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~3 .lut_mask = 16'hFCAA;
defparam \Mux31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N26
cycloneive_lcell_comb \ShiftRight0~30 (
// Equation(s):
// \ShiftRight0~30_combout  = (!Mux301 & ((Mux311 & ((alu_a_mux_output_1))) # (!Mux311 & (alu_a_mux_output_0))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_0),
	.datac(alu_a_mux_output_1),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftRight0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~30 .lut_mask = 16'h5044;
defparam \ShiftRight0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N2
cycloneive_lcell_comb \ShiftRight0~32 (
// Equation(s):
// \ShiftRight0~32_combout  = (!Mux291 & ((\ShiftRight0~30_combout ) # ((Mux301 & \ShiftRight0~31_combout ))))

	.dataa(Mux301),
	.datab(Mux291),
	.datac(\ShiftRight0~30_combout ),
	.datad(\ShiftRight0~31_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~32 .lut_mask = 16'h3230;
defparam \ShiftRight0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N16
cycloneive_lcell_comb \ShiftRight0~36 (
// Equation(s):
// \ShiftRight0~36_combout  = (!Mux281 & ((\ShiftRight0~32_combout ) # ((Mux291 & \ShiftRight0~35_combout ))))

	.dataa(Mux281),
	.datab(Mux291),
	.datac(\ShiftRight0~35_combout ),
	.datad(\ShiftRight0~32_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~36 .lut_mask = 16'h5540;
defparam \ShiftRight0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N6
cycloneive_lcell_comb \ShiftRight0~42 (
// Equation(s):
// \ShiftRight0~42_combout  = (!Mux271 & ((\ShiftRight0~36_combout ) # ((Mux281 & \ShiftRight0~41_combout ))))

	.dataa(Mux281),
	.datab(\ShiftRight0~41_combout ),
	.datac(Mux271),
	.datad(\ShiftRight0~36_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~42 .lut_mask = 16'h0F08;
defparam \ShiftRight0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N12
cycloneive_lcell_comb \ShiftRight0~50 (
// Equation(s):
// \ShiftRight0~50_combout  = (Mux301 & ((Mux311 & ((alu_a_mux_output_19))) # (!Mux311 & (alu_a_mux_output_18))))

	.dataa(Mux311),
	.datab(alu_a_mux_output_18),
	.datac(Mux301),
	.datad(alu_a_mux_output_19),
	.cin(gnd),
	.combout(\ShiftRight0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~50 .lut_mask = 16'hE040;
defparam \ShiftRight0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N28
cycloneive_lcell_comb \ShiftRight0~52 (
// Equation(s):
// \ShiftRight0~52_combout  = (Mux281 & (Mux291 & ((\ShiftRight0~45_combout )))) # (!Mux281 & (((\ShiftRight0~51_combout ))))

	.dataa(Mux281),
	.datab(Mux291),
	.datac(\ShiftRight0~51_combout ),
	.datad(\ShiftRight0~45_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~52 .lut_mask = 16'hD850;
defparam \ShiftRight0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N30
cycloneive_lcell_comb \Mux31~4 (
// Equation(s):
// \Mux31~4_combout  = (!\ShiftLeft0~11_combout  & ((\ShiftRight0~42_combout ) # ((\Mux31~3_combout  & \ShiftRight0~55_combout ))))

	.dataa(\Mux31~3_combout ),
	.datab(\ShiftLeft0~11_combout ),
	.datac(\ShiftRight0~55_combout ),
	.datad(\ShiftRight0~42_combout ),
	.cin(gnd),
	.combout(\Mux31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~4 .lut_mask = 16'h3320;
defparam \Mux31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N8
cycloneive_lcell_comb \Mux31~5 (
// Equation(s):
// \Mux31~5_combout  = (temp_ALUop_output_0 & (((\Mux31~4_combout )))) # (!temp_ALUop_output_0 & (\ShiftLeft0~17_combout  & ((!\Mux31~3_combout ))))

	.dataa(temp_ALUop_output_0),
	.datab(\ShiftLeft0~17_combout ),
	.datac(\Mux31~4_combout ),
	.datad(\Mux31~3_combout ),
	.cin(gnd),
	.combout(\Mux31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~5 .lut_mask = 16'hA0E4;
defparam \Mux31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N8
cycloneive_lcell_comb \ShiftRight0~63 (
// Equation(s):
// \ShiftRight0~63_combout  = (Mux301 & ((Mux311 & (alu_a_mux_output_17)) # (!Mux311 & ((alu_a_mux_output_16)))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_17),
	.datac(Mux311),
	.datad(alu_a_mux_output_16),
	.cin(gnd),
	.combout(\ShiftRight0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~63 .lut_mask = 16'h8A80;
defparam \ShiftRight0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N12
cycloneive_lcell_comb \ShiftRight0~69 (
// Equation(s):
// \ShiftRight0~69_combout  = (Mux311 & (((alu_a_mux_output_25) # (!Mux301)))) # (!Mux311 & (alu_a_mux_output_24 & (Mux301)))

	.dataa(Mux311),
	.datab(alu_a_mux_output_24),
	.datac(Mux301),
	.datad(alu_a_mux_output_25),
	.cin(gnd),
	.combout(\ShiftRight0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~69 .lut_mask = 16'hEA4A;
defparam \ShiftRight0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N14
cycloneive_lcell_comb \ShiftRight0~70 (
// Equation(s):
// \ShiftRight0~70_combout  = (Mux301 & (((\ShiftRight0~69_combout )))) # (!Mux301 & ((\ShiftRight0~69_combout  & (alu_a_mux_output_23)) # (!\ShiftRight0~69_combout  & ((alu_a_mux_output_22)))))

	.dataa(alu_a_mux_output_23),
	.datab(alu_a_mux_output_22),
	.datac(Mux301),
	.datad(\ShiftRight0~69_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~70 .lut_mask = 16'hFA0C;
defparam \ShiftRight0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N4
cycloneive_lcell_comb \ShiftLeft0~19 (
// Equation(s):
// \ShiftLeft0~19_combout  = (\ShiftRight0~59_combout  & ((\ShiftLeft0~18_combout ) # ((\Mux1~0_combout  & alu_a_mux_output_1))))

	.dataa(\Mux1~0_combout ),
	.datab(\ShiftRight0~59_combout ),
	.datac(alu_a_mux_output_1),
	.datad(\ShiftLeft0~18_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~19 .lut_mask = 16'hCC80;
defparam \ShiftLeft0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N6
cycloneive_lcell_comb \OUTPUT~0 (
// Equation(s):
// \OUTPUT~0_combout  = (alu_a_mux_output_2 & ((Mux29) # ((!Mux16 & alu_b_mux_output_2))))

	.dataa(alu_a_mux_output_2),
	.datab(Mux16),
	.datac(Mux29),
	.datad(alu_b_mux_output_2),
	.cin(gnd),
	.combout(\OUTPUT~0_combout ),
	.cout());
// synopsys translate_off
defparam \OUTPUT~0 .lut_mask = 16'hA2A0;
defparam \OUTPUT~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N16
cycloneive_lcell_comb \Mux29~6 (
// Equation(s):
// \Mux29~6_combout  = (\Mux29~5_combout  & ((\OUTPUT~0_combout ) # ((!\Mux29~4_combout )))) # (!\Mux29~5_combout  & (((\ShiftLeft0~19_combout  & \Mux29~4_combout ))))

	.dataa(\OUTPUT~0_combout ),
	.datab(\Mux29~5_combout ),
	.datac(\ShiftLeft0~19_combout ),
	.datad(\Mux29~4_combout ),
	.cin(gnd),
	.combout(\Mux29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~6 .lut_mask = 16'hB8CC;
defparam \Mux29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N22
cycloneive_lcell_comb \OUTPUT~1 (
// Equation(s):
// \OUTPUT~1_combout  = (alu_a_mux_output_31 & ((Mux28) # ((!Mux16 & alu_b_mux_output_3))))

	.dataa(alu_a_mux_output_31),
	.datab(Mux16),
	.datac(Mux28),
	.datad(alu_b_mux_output_3),
	.cin(gnd),
	.combout(\OUTPUT~1_combout ),
	.cout());
// synopsys translate_off
defparam \OUTPUT~1 .lut_mask = 16'hA2A0;
defparam \OUTPUT~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N4
cycloneive_lcell_comb \Mux26~2 (
// Equation(s):
// \Mux26~2_combout  = (!Mux281 & (\Mux19~0_combout  & \ShiftLeft0~25_combout ))

	.dataa(Mux281),
	.datab(gnd),
	.datac(\Mux19~0_combout ),
	.datad(\ShiftLeft0~25_combout ),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~2 .lut_mask = 16'h5000;
defparam \Mux26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N14
cycloneive_lcell_comb \ShiftLeft0~27 (
// Equation(s):
// \ShiftLeft0~27_combout  = (Mux301 & (((alu_a_mux_output_1)))) # (!Mux301 & ((alu_a_mux_output_3) # ((alu_a_mux_output_32))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_3),
	.datac(alu_a_mux_output_32),
	.datad(alu_a_mux_output_1),
	.cin(gnd),
	.combout(\ShiftLeft0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~27 .lut_mask = 16'hFE54;
defparam \ShiftLeft0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N10
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (\Mux27~3_combout  & (((\ShiftRight0~96_combout ) # (\Mux27~2_combout )))) # (!\Mux27~3_combout  & (\ShiftRight0~75_combout  & ((!\Mux27~2_combout ))))

	.dataa(\Mux27~3_combout ),
	.datab(\ShiftRight0~75_combout ),
	.datac(\ShiftRight0~96_combout ),
	.datad(\Mux27~2_combout ),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hAAE4;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N26
cycloneive_lcell_comb \ShiftLeft0~38 (
// Equation(s):
// \ShiftLeft0~38_combout  = (Mux301 & ((alu_a_mux_output_7))) # (!Mux301 & (alu_a_mux_output_9))

	.dataa(Mux301),
	.datab(gnd),
	.datac(alu_a_mux_output_9),
	.datad(alu_a_mux_output_7),
	.cin(gnd),
	.combout(\ShiftLeft0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~38 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N0
cycloneive_lcell_comb \ShiftLeft0~42 (
// Equation(s):
// \ShiftLeft0~42_combout  = (Mux311 & ((Mux301 & ((alu_a_mux_output_5))) # (!Mux301 & (alu_a_mux_output_7))))

	.dataa(Mux311),
	.datab(Mux301),
	.datac(alu_a_mux_output_7),
	.datad(alu_a_mux_output_5),
	.cin(gnd),
	.combout(\ShiftLeft0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~42 .lut_mask = 16'hA820;
defparam \ShiftLeft0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N2
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (!\ShiftLeft0~26_combout  & (\ShiftLeft0~50_combout  & (!\ShiftLeft0~10_combout  & !Mux271)))

	.dataa(\ShiftLeft0~26_combout ),
	.datab(\ShiftLeft0~50_combout ),
	.datac(\ShiftLeft0~10_combout ),
	.datad(Mux271),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'h0004;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N10
cycloneive_lcell_comb \ShiftRight0~106 (
// Equation(s):
// \ShiftRight0~106_combout  = (!Mux301 & (!Mux281 & (Mux291 & \ShiftRight0~44_combout )))

	.dataa(Mux301),
	.datab(Mux281),
	.datac(Mux291),
	.datad(\ShiftRight0~44_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~106_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~106 .lut_mask = 16'h1000;
defparam \ShiftRight0~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N12
cycloneive_lcell_comb \Mux19~8 (
// Equation(s):
// \Mux19~8_combout  = (!Mux271 & (!\ShiftLeft0~26_combout  & (!\ShiftLeft0~10_combout  & \ShiftLeft0~61_combout )))

	.dataa(Mux271),
	.datab(\ShiftLeft0~26_combout ),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\ShiftLeft0~61_combout ),
	.cin(gnd),
	.combout(\Mux19~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~8 .lut_mask = 16'h0100;
defparam \Mux19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N28
cycloneive_lcell_comb \ShiftLeft0~75 (
// Equation(s):
// \ShiftLeft0~75_combout  = (!Mux311 & ((Mux301 & (alu_a_mux_output_17)) # (!Mux301 & ((alu_a_mux_output_19)))))

	.dataa(alu_a_mux_output_17),
	.datab(Mux301),
	.datac(Mux311),
	.datad(alu_a_mux_output_19),
	.cin(gnd),
	.combout(\ShiftLeft0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~75 .lut_mask = 16'h0B08;
defparam \ShiftLeft0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N4
cycloneive_lcell_comb \Mux12~4 (
// Equation(s):
// \Mux12~4_combout  = (\ShiftRight0~59_combout  & (!\ShiftLeft0~10_combout  & (!\ShiftLeft0~26_combout  & \ShiftLeft0~30_combout )))

	.dataa(\ShiftRight0~59_combout ),
	.datab(\ShiftLeft0~10_combout ),
	.datac(\ShiftLeft0~26_combout ),
	.datad(\ShiftLeft0~30_combout ),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~4 .lut_mask = 16'h0200;
defparam \Mux12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N10
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (\ShiftLeft0~104_combout  & (!\ShiftLeft0~26_combout  & (!\ShiftLeft0~10_combout  & \ShiftRight0~59_combout )))

	.dataa(\ShiftLeft0~104_combout ),
	.datab(\ShiftLeft0~26_combout ),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\ShiftRight0~59_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'h0200;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N26
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (!temp_ALUop_output_1 & ((\Mux19~0_combout ) # (!temp_ALUop_output_0)))

	.dataa(temp_ALUop_output_0),
	.datab(temp_ALUop_output_1),
	.datac(\Mux19~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'h3131;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N4
cycloneive_lcell_comb \ShiftLeft0~99 (
// Equation(s):
// \ShiftLeft0~99_combout  = (Mux301 & ((Mux311 & ((alu_a_mux_output_24))) # (!Mux311 & (alu_a_mux_output_25))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_25),
	.datac(Mux311),
	.datad(alu_a_mux_output_24),
	.cin(gnd),
	.combout(\ShiftLeft0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~99 .lut_mask = 16'hA808;
defparam \ShiftLeft0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N10
cycloneive_lcell_comb \ShiftLeft0~100 (
// Equation(s):
// \ShiftLeft0~100_combout  = (Mux311 & (alu_a_mux_output_26)) # (!Mux311 & ((alu_a_mux_output_27)))

	.dataa(gnd),
	.datab(alu_a_mux_output_26),
	.datac(Mux311),
	.datad(alu_a_mux_output_27),
	.cin(gnd),
	.combout(\ShiftLeft0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~100 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N0
cycloneive_lcell_comb \ShiftLeft0~101 (
// Equation(s):
// \ShiftLeft0~101_combout  = (\ShiftLeft0~99_combout ) # ((!Mux301 & \ShiftLeft0~100_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~99_combout ),
	.datac(Mux301),
	.datad(\ShiftLeft0~100_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~101 .lut_mask = 16'hCFCC;
defparam \ShiftLeft0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N6
cycloneive_lcell_comb \Mux4~2 (
// Equation(s):
// \Mux4~2_combout  = (\Mux27~3_combout  & (((\Mux27~2_combout ) # (\ShiftLeft0~76_combout )))) # (!\Mux27~3_combout  & (\ShiftLeft0~101_combout  & (!\Mux27~2_combout )))

	.dataa(\ShiftLeft0~101_combout ),
	.datab(\Mux27~3_combout ),
	.datac(\Mux27~2_combout ),
	.datad(\ShiftLeft0~76_combout ),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~2 .lut_mask = 16'hCEC2;
defparam \Mux4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N12
cycloneive_lcell_comb \ShiftLeft0~103 (
// Equation(s):
// \ShiftLeft0~103_combout  = (Mux311 & ((alu_a_mux_output_27))) # (!Mux311 & (alu_a_mux_output_28))

	.dataa(gnd),
	.datab(alu_a_mux_output_28),
	.datac(Mux311),
	.datad(alu_a_mux_output_27),
	.cin(gnd),
	.combout(\ShiftLeft0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~103 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N4
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (\ShiftRight0~59_combout  & (\ShiftLeft0~103_combout  & ((!\Mux29~0_combout )))) # (!\ShiftRight0~59_combout  & (((\ShiftLeft0~95_combout ) # (\Mux29~0_combout ))))

	.dataa(\ShiftRight0~59_combout ),
	.datab(\ShiftLeft0~103_combout ),
	.datac(\ShiftLeft0~95_combout ),
	.datad(\Mux29~0_combout ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'h55D8;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N26
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (\Mux3~0_combout  & (((\ShiftLeft0~82_combout ) # (!\Mux29~0_combout )))) # (!\Mux3~0_combout  & (\ShiftLeft0~97_combout  & ((\Mux29~0_combout ))))

	.dataa(\ShiftLeft0~97_combout ),
	.datab(\ShiftLeft0~82_combout ),
	.datac(\Mux3~0_combout ),
	.datad(\Mux29~0_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hCAF0;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N14
cycloneive_lcell_comb \OUTPUT~3 (
// Equation(s):
// \OUTPUT~3_combout  = (alu_a_mux_output_28 & Mux3)

	.dataa(gnd),
	.datab(alu_a_mux_output_28),
	.datac(gnd),
	.datad(Mux3),
	.cin(gnd),
	.combout(\OUTPUT~3_combout ),
	.cout());
// synopsys translate_off
defparam \OUTPUT~3 .lut_mask = 16'hCC00;
defparam \OUTPUT~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N18
cycloneive_lcell_comb \Mux10~6 (
// Equation(s):
// \Mux10~6_combout  = (temp_ALUop_output_2 & (((Mux102)))) # (!temp_ALUop_output_2 & ((temp_ALUop_output_1 & (Mux101)) # (!temp_ALUop_output_1 & ((Mux102)))))

	.dataa(Mux101),
	.datab(temp_ALUop_output_2),
	.datac(Mux102),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Mux10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~6 .lut_mask = 16'hE2F0;
defparam \Mux10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N20
cycloneive_lcell_comb \Equal0~15 (
// Equation(s):
// \Equal0~15_combout  = (temp_ALUop_output_2 & (\Equal0~23_combout )) # (!temp_ALUop_output_2 & (((!Mux151 & !Mux01))))

	.dataa(temp_ALUop_output_2),
	.datab(\Equal0~23_combout ),
	.datac(Mux151),
	.datad(Mux01),
	.cin(gnd),
	.combout(\Equal0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~15 .lut_mask = 16'h888D;
defparam \Equal0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N22
cycloneive_lcell_comb \Equal0~16 (
// Equation(s):
// \Equal0~16_combout  = (temp_ALUop_output_1 & (\Equal0~15_combout  & ((!Mux152) # (!temp_ALUop_output_2)))) # (!temp_ALUop_output_1 & (((!Mux152))))

	.dataa(temp_ALUop_output_2),
	.datab(temp_ALUop_output_1),
	.datac(Mux152),
	.datad(\Equal0~15_combout ),
	.cin(gnd),
	.combout(\Equal0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~16 .lut_mask = 16'h4F03;
defparam \Equal0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N10
cycloneive_lcell_comb \Equal0~18 (
// Equation(s):
// \Equal0~18_combout  = (temp_ALUop_output_2 & (\Equal0~17_combout )) # (!temp_ALUop_output_2 & (((Mux151) # (Mux01))))

	.dataa(temp_ALUop_output_2),
	.datab(\Equal0~17_combout ),
	.datac(Mux151),
	.datad(Mux01),
	.cin(gnd),
	.combout(\Equal0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~18 .lut_mask = 16'hDDD8;
defparam \Equal0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N24
cycloneive_lcell_comb \Add0~105 (
// Equation(s):
// \Add0~105_combout  = (!Mux30 & ((temp_ALUsrc_output_1 $ (temp_ALUsrc_output_0)) # (!alu_b_mux_output_1)))

	.dataa(temp_ALUsrc_output_1),
	.datab(temp_ALUsrc_output_0),
	.datac(Mux30),
	.datad(alu_b_mux_output_1),
	.cin(gnd),
	.combout(\Add0~105_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~105 .lut_mask = 16'h060F;
defparam \Add0~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N30
cycloneive_lcell_comb \Mux2~15 (
// Equation(s):
// \Mux2~15_combout  = (temp_ALUop_output_1) # ((!temp_ALUop_output_2 & ((temp_ALUop_output_0) # (!\ShiftLeft0~11_combout ))))

	.dataa(temp_ALUop_output_2),
	.datab(temp_ALUop_output_1),
	.datac(\ShiftLeft0~11_combout ),
	.datad(temp_ALUop_output_0),
	.cin(gnd),
	.combout(\Mux2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~15 .lut_mask = 16'hDDCD;
defparam \Mux2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N20
cycloneive_lcell_comb \Mux30~4 (
// Equation(s):
// Mux302 = (!temp_ALUop_output_3 & ((temp_ALUop_output_2 & ((\Mux30~1_combout ))) # (!temp_ALUop_output_2 & (\Mux30~3_combout ))))

	.dataa(\Mux30~3_combout ),
	.datab(\Mux30~1_combout ),
	.datac(temp_ALUop_output_2),
	.datad(temp_ALUop_output_3),
	.cin(gnd),
	.combout(Mux302),
	.cout());
// synopsys translate_off
defparam \Mux30~4 .lut_mask = 16'h00CA;
defparam \Mux30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N8
cycloneive_lcell_comb \Mux31~9 (
// Equation(s):
// Mux312 = (\Mux31~8_combout  & ((temp_ALUop_output_0) # ((\LessThan0~62_combout ) # (!temp_ALUop_output_3))))

	.dataa(temp_ALUop_output_0),
	.datab(temp_ALUop_output_3),
	.datac(\LessThan0~62_combout ),
	.datad(\Mux31~8_combout ),
	.cin(gnd),
	.combout(Mux312),
	.cout());
// synopsys translate_off
defparam \Mux31~9 .lut_mask = 16'hFB00;
defparam \Mux31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N10
cycloneive_lcell_comb \Mux29~12 (
// Equation(s):
// Mux292 = (\Mux29~11_combout  & (((alu_a_mux_output_2) # (Mux291)))) # (!\Mux29~11_combout  & (\Mux29~10_combout ))

	.dataa(\Mux29~11_combout ),
	.datab(\Mux29~10_combout ),
	.datac(alu_a_mux_output_2),
	.datad(Mux291),
	.cin(gnd),
	.combout(Mux292),
	.cout());
// synopsys translate_off
defparam \Mux29~12 .lut_mask = 16'hEEE4;
defparam \Mux29~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N24
cycloneive_lcell_comb \Mux28~6 (
// Equation(s):
// Mux282 = (\Mux29~11_combout  & (((alu_a_mux_output_31) # (Mux281)))) # (!\Mux29~11_combout  & (\Mux28~5_combout ))

	.dataa(\Mux28~5_combout ),
	.datab(alu_a_mux_output_31),
	.datac(Mux281),
	.datad(\Mux29~11_combout ),
	.cin(gnd),
	.combout(Mux282),
	.cout());
// synopsys translate_off
defparam \Mux28~6 .lut_mask = 16'hFCAA;
defparam \Mux28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N12
cycloneive_lcell_comb \Mux26~6 (
// Equation(s):
// Mux261 = (\Mux26~5_combout  & ((\Add0~23_combout ) # ((!\Mux19~1_combout )))) # (!\Mux26~5_combout  & (((\Mux26~4_combout  & \Mux19~1_combout ))))

	.dataa(\Mux26~5_combout ),
	.datab(\Add0~23_combout ),
	.datac(\Mux26~4_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(Mux261),
	.cout());
// synopsys translate_off
defparam \Mux26~6 .lut_mask = 16'hD8AA;
defparam \Mux26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N28
cycloneive_lcell_comb \Mux27~11 (
// Equation(s):
// Mux272 = (\Mux27~10_combout  & (((\Add0~21_combout )) # (!\Mux19~1_combout ))) # (!\Mux27~10_combout  & (\Mux19~1_combout  & ((\Mux27~9_combout ))))

	.dataa(\Mux27~10_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Add0~21_combout ),
	.datad(\Mux27~9_combout ),
	.cin(gnd),
	.combout(Mux272),
	.cout());
// synopsys translate_off
defparam \Mux27~11 .lut_mask = 16'hE6A2;
defparam \Mux27~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N20
cycloneive_lcell_comb \Mux24~6 (
// Equation(s):
// Mux241 = (\Mux24~5_combout  & (((\Add0~31_combout )) # (!\Mux19~1_combout ))) # (!\Mux24~5_combout  & (\Mux19~1_combout  & (\Mux24~4_combout )))

	.dataa(\Mux24~5_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Mux24~4_combout ),
	.datad(\Add0~31_combout ),
	.cin(gnd),
	.combout(Mux241),
	.cout());
// synopsys translate_off
defparam \Mux24~6 .lut_mask = 16'hEA62;
defparam \Mux24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N10
cycloneive_lcell_comb \Mux25~6 (
// Equation(s):
// Mux251 = (\Mux19~1_combout  & ((\Mux25~5_combout  & (\Add0~29_combout )) # (!\Mux25~5_combout  & ((\Mux25~4_combout ))))) # (!\Mux19~1_combout  & (((\Mux25~5_combout ))))

	.dataa(\Add0~29_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Mux25~5_combout ),
	.datad(\Mux25~4_combout ),
	.cin(gnd),
	.combout(Mux251),
	.cout());
// synopsys translate_off
defparam \Mux25~6 .lut_mask = 16'hBCB0;
defparam \Mux25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N20
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// Mux221 = (alu_a_mux_output_9 & ((temp_ALUop_output_0) # (Mux22))) # (!alu_a_mux_output_9 & (temp_ALUop_output_0 & Mux22))

	.dataa(gnd),
	.datab(alu_a_mux_output_9),
	.datac(temp_ALUop_output_0),
	.datad(Mux22),
	.cin(gnd),
	.combout(Mux221),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hFCC0;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N22
cycloneive_lcell_comb \Mux22~5 (
// Equation(s):
// Mux222 = (\Mux19~1_combout  & ((\Mux22~4_combout  & ((\Add0~37_combout ))) # (!\Mux22~4_combout  & (\Mux22~3_combout )))) # (!\Mux19~1_combout  & (((\Mux22~4_combout ))))

	.dataa(\Mux22~3_combout ),
	.datab(\Add0~37_combout ),
	.datac(\Mux19~1_combout ),
	.datad(\Mux22~4_combout ),
	.cin(gnd),
	.combout(Mux222),
	.cout());
// synopsys translate_off
defparam \Mux22~5 .lut_mask = 16'hCFA0;
defparam \Mux22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N18
cycloneive_lcell_comb \Mux19~6 (
// Equation(s):
// Mux191 = (!temp_ALUop_output_2 & temp_ALUop_output_1)

	.dataa(temp_ALUop_output_2),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(Mux191),
	.cout());
// synopsys translate_off
defparam \Mux19~6 .lut_mask = 16'h5500;
defparam \Mux19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N12
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// Mux231 = (Mux191 & ((alu_a_mux_output_8 & ((Mux23) # (temp_ALUop_output_0))) # (!alu_a_mux_output_8 & (Mux23 & temp_ALUop_output_0))))

	.dataa(alu_a_mux_output_8),
	.datab(Mux191),
	.datac(Mux23),
	.datad(temp_ALUop_output_0),
	.cin(gnd),
	.combout(Mux231),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hC880;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N4
cycloneive_lcell_comb \Mux23~5 (
// Equation(s):
// Mux232 = (\Mux19~1_combout  & ((\Mux23~4_combout  & (\Add0~35_combout )) # (!\Mux23~4_combout  & ((\Mux23~3_combout ))))) # (!\Mux19~1_combout  & (((\Mux23~4_combout ))))

	.dataa(\Add0~35_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Mux23~4_combout ),
	.datad(\Mux23~3_combout ),
	.cin(gnd),
	.combout(Mux232),
	.cout());
// synopsys translate_off
defparam \Mux23~5 .lut_mask = 16'hBCB0;
defparam \Mux23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N22
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// Mux201 = (temp_ALUop_output_0 & ((alu_a_mux_output_11) # (Mux20))) # (!temp_ALUop_output_0 & (alu_a_mux_output_11 & Mux20))

	.dataa(temp_ALUop_output_0),
	.datab(alu_a_mux_output_11),
	.datac(Mux20),
	.datad(gnd),
	.cin(gnd),
	.combout(Mux201),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hE8E8;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y43_N10
cycloneive_lcell_comb \Mux20~5 (
// Equation(s):
// Mux202 = (\Mux20~4_combout  & (((\Add0~43_combout )) # (!\Mux19~1_combout ))) # (!\Mux20~4_combout  & (\Mux19~1_combout  & ((\Mux20~3_combout ))))

	.dataa(\Mux20~4_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Add0~43_combout ),
	.datad(\Mux20~3_combout ),
	.cin(gnd),
	.combout(Mux202),
	.cout());
// synopsys translate_off
defparam \Mux20~5 .lut_mask = 16'hE6A2;
defparam \Mux20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N4
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// Mux211 = (temp_ALUop_output_0 & ((alu_a_mux_output_10) # (Mux21))) # (!temp_ALUop_output_0 & (alu_a_mux_output_10 & Mux21))

	.dataa(temp_ALUop_output_0),
	.datab(alu_a_mux_output_10),
	.datac(gnd),
	.datad(Mux21),
	.cin(gnd),
	.combout(Mux211),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hEE88;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y43_N26
cycloneive_lcell_comb \Mux21~5 (
// Equation(s):
// Mux212 = (\Mux21~4_combout  & (((\Add0~41_combout ) # (!\Mux19~1_combout )))) # (!\Mux21~4_combout  & (\Mux21~3_combout  & (\Mux19~1_combout )))

	.dataa(\Mux21~3_combout ),
	.datab(\Mux21~4_combout ),
	.datac(\Mux19~1_combout ),
	.datad(\Add0~41_combout ),
	.cin(gnd),
	.combout(Mux212),
	.cout());
// synopsys translate_off
defparam \Mux21~5 .lut_mask = 16'hEC2C;
defparam \Mux21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N24
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// Mux181 = (temp_ALUop_output_0 & ((alu_a_mux_output_13) # (Mux18))) # (!temp_ALUop_output_0 & (alu_a_mux_output_13 & Mux18))

	.dataa(temp_ALUop_output_0),
	.datab(alu_a_mux_output_13),
	.datac(Mux18),
	.datad(gnd),
	.cin(gnd),
	.combout(Mux181),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hE8E8;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N16
cycloneive_lcell_comb \Mux18~5 (
// Equation(s):
// Mux182 = (\Mux19~1_combout  & ((\Mux18~4_combout  & (\Add0~49_combout )) # (!\Mux18~4_combout  & ((\Mux18~3_combout ))))) # (!\Mux19~1_combout  & (((\Mux18~4_combout ))))

	.dataa(\Add0~49_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Mux18~3_combout ),
	.datad(\Mux18~4_combout ),
	.cin(gnd),
	.combout(Mux182),
	.cout());
// synopsys translate_off
defparam \Mux18~5 .lut_mask = 16'hBBC0;
defparam \Mux18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N6
cycloneive_lcell_comb \Mux19~7 (
// Equation(s):
// Mux192 = (Mux19 & ((temp_ALUop_output_0) # (alu_a_mux_output_12))) # (!Mux19 & (temp_ALUop_output_0 & alu_a_mux_output_12))

	.dataa(gnd),
	.datab(Mux19),
	.datac(temp_ALUop_output_0),
	.datad(alu_a_mux_output_12),
	.cin(gnd),
	.combout(Mux192),
	.cout());
// synopsys translate_off
defparam \Mux19~7 .lut_mask = 16'hFCC0;
defparam \Mux19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N14
cycloneive_lcell_comb \Mux19~12 (
// Equation(s):
// Mux193 = (\Mux19~11_combout  & ((\Add0~47_combout ) # ((!\Mux19~1_combout )))) # (!\Mux19~11_combout  & (((\Mux19~1_combout  & \Mux19~10_combout ))))

	.dataa(\Add0~47_combout ),
	.datab(\Mux19~11_combout ),
	.datac(\Mux19~1_combout ),
	.datad(\Mux19~10_combout ),
	.cin(gnd),
	.combout(Mux193),
	.cout());
// synopsys translate_off
defparam \Mux19~12 .lut_mask = 16'hBC8C;
defparam \Mux19~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N22
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// Mux162 = (Mux161 & ((alu_a_mux_output_15) # (temp_ALUop_output_0))) # (!Mux161 & (alu_a_mux_output_15 & temp_ALUop_output_0))

	.dataa(Mux161),
	.datab(alu_a_mux_output_15),
	.datac(temp_ALUop_output_0),
	.datad(gnd),
	.cin(gnd),
	.combout(Mux162),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hE8E8;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N14
cycloneive_lcell_comb \Mux16~5 (
// Equation(s):
// Mux163 = (\Mux16~4_combout  & ((\Add0~55_combout ) # ((!\Mux19~1_combout )))) # (!\Mux16~4_combout  & (((\Mux16~3_combout  & \Mux19~1_combout ))))

	.dataa(\Mux16~4_combout ),
	.datab(\Add0~55_combout ),
	.datac(\Mux16~3_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(Mux163),
	.cout());
// synopsys translate_off
defparam \Mux16~5 .lut_mask = 16'hD8AA;
defparam \Mux16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N0
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// Mux172 = (Mux171 & ((alu_a_mux_output_14) # (temp_ALUop_output_0))) # (!Mux171 & (alu_a_mux_output_14 & temp_ALUop_output_0))

	.dataa(Mux171),
	.datab(alu_a_mux_output_14),
	.datac(gnd),
	.datad(temp_ALUop_output_0),
	.cin(gnd),
	.combout(Mux172),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hEE88;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N0
cycloneive_lcell_comb \Mux17~5 (
// Equation(s):
// Mux173 = (\Mux19~1_combout  & ((\Mux17~4_combout  & (\Add0~53_combout )) # (!\Mux17~4_combout  & ((\Mux17~3_combout ))))) # (!\Mux19~1_combout  & (((\Mux17~4_combout ))))

	.dataa(\Add0~53_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Mux17~4_combout ),
	.datad(\Mux17~3_combout ),
	.cin(gnd),
	.combout(Mux173),
	.cout());
// synopsys translate_off
defparam \Mux17~5 .lut_mask = 16'hBCB0;
defparam \Mux17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N0
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// Mux141 = (temp_ALUop_output_0 & ((Mux14) # (alu_a_mux_output_17))) # (!temp_ALUop_output_0 & (Mux14 & alu_a_mux_output_17))

	.dataa(gnd),
	.datab(temp_ALUop_output_0),
	.datac(Mux14),
	.datad(alu_a_mux_output_17),
	.cin(gnd),
	.combout(Mux141),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hFCC0;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N20
cycloneive_lcell_comb \Mux14~4 (
// Equation(s):
// Mux142 = (\Mux19~1_combout  & ((\Mux14~3_combout  & ((\Add0~61_combout ))) # (!\Mux14~3_combout  & (\Mux14~2_combout )))) # (!\Mux19~1_combout  & (((\Mux14~3_combout ))))

	.dataa(\Mux19~1_combout ),
	.datab(\Mux14~2_combout ),
	.datac(\Mux14~3_combout ),
	.datad(\Add0~61_combout ),
	.cin(gnd),
	.combout(Mux142),
	.cout());
// synopsys translate_off
defparam \Mux14~4 .lut_mask = 16'hF858;
defparam \Mux14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N4
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// Mux151 = (Mux15 & ((temp_ALUop_output_0) # (alu_a_mux_output_16))) # (!Mux15 & (temp_ALUop_output_0 & alu_a_mux_output_16))

	.dataa(gnd),
	.datab(Mux15),
	.datac(temp_ALUop_output_0),
	.datad(alu_a_mux_output_16),
	.cin(gnd),
	.combout(Mux151),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hFCC0;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N8
cycloneive_lcell_comb \Mux15~4 (
// Equation(s):
// Mux152 = (\Mux19~1_combout  & ((\Mux15~3_combout  & (\Add0~59_combout )) # (!\Mux15~3_combout  & ((\Mux15~2_combout ))))) # (!\Mux19~1_combout  & (((\Mux15~3_combout ))))

	.dataa(\Add0~59_combout ),
	.datab(\Mux15~2_combout ),
	.datac(\Mux19~1_combout ),
	.datad(\Mux15~3_combout ),
	.cin(gnd),
	.combout(Mux152),
	.cout());
// synopsys translate_off
defparam \Mux15~4 .lut_mask = 16'hAFC0;
defparam \Mux15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N22
cycloneive_lcell_comb \Mux12~3 (
// Equation(s):
// Mux121 = (Mux12 & ((temp_ALUop_output_0) # (alu_a_mux_output_19))) # (!Mux12 & (temp_ALUop_output_0 & alu_a_mux_output_19))

	.dataa(gnd),
	.datab(Mux12),
	.datac(temp_ALUop_output_0),
	.datad(alu_a_mux_output_19),
	.cin(gnd),
	.combout(Mux121),
	.cout());
// synopsys translate_off
defparam \Mux12~3 .lut_mask = 16'hFCC0;
defparam \Mux12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N30
cycloneive_lcell_comb \Mux12~8 (
// Equation(s):
// Mux122 = (\Mux19~1_combout  & ((\Mux12~7_combout  & (\Add0~67_combout )) # (!\Mux12~7_combout  & ((\Mux12~6_combout ))))) # (!\Mux19~1_combout  & (((\Mux12~7_combout ))))

	.dataa(\Add0~67_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Mux12~6_combout ),
	.datad(\Mux12~7_combout ),
	.cin(gnd),
	.combout(Mux122),
	.cout());
// synopsys translate_off
defparam \Mux12~8 .lut_mask = 16'hBBC0;
defparam \Mux12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N10
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// Mux131 = (Mux13 & ((alu_a_mux_output_18) # (temp_ALUop_output_0))) # (!Mux13 & (alu_a_mux_output_18 & temp_ALUop_output_0))

	.dataa(gnd),
	.datab(Mux13),
	.datac(alu_a_mux_output_18),
	.datad(temp_ALUop_output_0),
	.cin(gnd),
	.combout(Mux131),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hFCC0;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N18
cycloneive_lcell_comb \Mux13~5 (
// Equation(s):
// Mux132 = (\Mux19~1_combout  & ((\Mux13~4_combout  & ((\Add0~65_combout ))) # (!\Mux13~4_combout  & (\Mux13~3_combout )))) # (!\Mux19~1_combout  & (\Mux13~4_combout ))

	.dataa(\Mux19~1_combout ),
	.datab(\Mux13~4_combout ),
	.datac(\Mux13~3_combout ),
	.datad(\Add0~65_combout ),
	.cin(gnd),
	.combout(Mux132),
	.cout());
// synopsys translate_off
defparam \Mux13~5 .lut_mask = 16'hEC64;
defparam \Mux13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N18
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// Mux111 = (alu_a_mux_output_20 & ((temp_ALUop_output_0) # (Mux11))) # (!alu_a_mux_output_20 & (temp_ALUop_output_0 & Mux11))

	.dataa(gnd),
	.datab(alu_a_mux_output_20),
	.datac(temp_ALUop_output_0),
	.datad(Mux11),
	.cin(gnd),
	.combout(Mux111),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hFCC0;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y43_N8
cycloneive_lcell_comb \Mux11~5 (
// Equation(s):
// Mux112 = (\Mux19~1_combout  & ((\Mux11~4_combout  & ((\Add0~70_combout ))) # (!\Mux11~4_combout  & (\Mux11~3_combout )))) # (!\Mux19~1_combout  & (((\Mux11~4_combout ))))

	.dataa(\Mux11~3_combout ),
	.datab(\Add0~70_combout ),
	.datac(\Mux19~1_combout ),
	.datad(\Mux11~4_combout ),
	.cin(gnd),
	.combout(Mux112),
	.cout());
// synopsys translate_off
defparam \Mux11~5 .lut_mask = 16'hCFA0;
defparam \Mux11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N2
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// Mux101 = (temp_ALUop_output_0 & ((alu_a_mux_output_21) # (Mux10))) # (!temp_ALUop_output_0 & (alu_a_mux_output_21 & Mux10))

	.dataa(gnd),
	.datab(temp_ALUop_output_0),
	.datac(alu_a_mux_output_21),
	.datad(Mux10),
	.cin(gnd),
	.combout(Mux101),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hFCC0;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N18
cycloneive_lcell_comb \Mux10~5 (
// Equation(s):
// Mux102 = (\Mux19~1_combout  & ((\Mux10~4_combout  & (\Add0~73_combout )) # (!\Mux10~4_combout  & ((\Mux10~3_combout ))))) # (!\Mux19~1_combout  & (((\Mux10~4_combout ))))

	.dataa(\Add0~73_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Mux10~3_combout ),
	.datad(\Mux10~4_combout ),
	.cin(gnd),
	.combout(Mux102),
	.cout());
// synopsys translate_off
defparam \Mux10~5 .lut_mask = 16'hBBC0;
defparam \Mux10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N18
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// Mux81 = (Mux8 & ((temp_ALUop_output_0) # (alu_a_mux_output_23))) # (!Mux8 & (temp_ALUop_output_0 & alu_a_mux_output_23))

	.dataa(gnd),
	.datab(Mux8),
	.datac(temp_ALUop_output_0),
	.datad(alu_a_mux_output_23),
	.cin(gnd),
	.combout(Mux81),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hFCC0;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N26
cycloneive_lcell_comb \Mux8~5 (
// Equation(s):
// Mux82 = (\Mux8~4_combout  & (((\Add0~79_combout )) # (!\Mux19~1_combout ))) # (!\Mux8~4_combout  & (\Mux19~1_combout  & (\Mux8~3_combout )))

	.dataa(\Mux8~4_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Mux8~3_combout ),
	.datad(\Add0~79_combout ),
	.cin(gnd),
	.combout(Mux82),
	.cout());
// synopsys translate_off
defparam \Mux8~5 .lut_mask = 16'hEA62;
defparam \Mux8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N2
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// Mux91 = (Mux191 & ((Mux9 & ((alu_a_mux_output_22) # (temp_ALUop_output_0))) # (!Mux9 & (alu_a_mux_output_22 & temp_ALUop_output_0))))

	.dataa(Mux9),
	.datab(alu_a_mux_output_22),
	.datac(temp_ALUop_output_0),
	.datad(Mux191),
	.cin(gnd),
	.combout(Mux91),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hE800;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N10
cycloneive_lcell_comb \Mux9~5 (
// Equation(s):
// Mux92 = (\Mux9~4_combout  & (((\Add0~77_combout ) # (!\Mux19~1_combout )))) # (!\Mux9~4_combout  & (\Mux9~3_combout  & ((\Mux19~1_combout ))))

	.dataa(\Mux9~4_combout ),
	.datab(\Mux9~3_combout ),
	.datac(\Add0~77_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(Mux92),
	.cout());
// synopsys translate_off
defparam \Mux9~5 .lut_mask = 16'hE4AA;
defparam \Mux9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N24
cycloneive_lcell_comb \Mux6~7 (
// Equation(s):
// Mux61 = (\Mux6~6_combout  & (((\Add0~85_combout )) # (!\Mux19~1_combout ))) # (!\Mux6~6_combout  & (\Mux19~1_combout  & (\Mux6~5_combout )))

	.dataa(\Mux6~6_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Mux6~5_combout ),
	.datad(\Add0~85_combout ),
	.cin(gnd),
	.combout(Mux61),
	.cout());
// synopsys translate_off
defparam \Mux6~7 .lut_mask = 16'hEA62;
defparam \Mux6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y43_N16
cycloneive_lcell_comb \Mux4~7 (
// Equation(s):
// Mux41 = (\Mux19~1_combout  & ((\Mux4~6_combout  & ((\Add0~91_combout ))) # (!\Mux4~6_combout  & (\Mux4~5_combout )))) # (!\Mux19~1_combout  & (((\Mux4~6_combout ))))

	.dataa(\Mux4~5_combout ),
	.datab(\Mux19~1_combout ),
	.datac(\Add0~91_combout ),
	.datad(\Mux4~6_combout ),
	.cin(gnd),
	.combout(Mux41),
	.cout());
// synopsys translate_off
defparam \Mux4~7 .lut_mask = 16'hF388;
defparam \Mux4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N30
cycloneive_lcell_comb \Mux2~14 (
// Equation(s):
// Mux210 = (\Mux29~11_combout  & (((\Mux2~13_combout )))) # (!\Mux29~11_combout  & ((\Add0~97_combout  & ((\Mux2~13_combout ))) # (!\Add0~97_combout  & (\Mux2~10_combout ))))

	.dataa(\Mux2~10_combout ),
	.datab(\Mux2~13_combout ),
	.datac(\Mux29~11_combout ),
	.datad(\Add0~97_combout ),
	.cin(gnd),
	.combout(Mux210),
	.cout());
// synopsys translate_off
defparam \Mux2~14 .lut_mask = 16'hCCCA;
defparam \Mux2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N2
cycloneive_lcell_comb \Mux3~9 (
// Equation(s):
// Mux32 = (\Add0~95_combout  & (((\Mux3~8_combout )))) # (!\Add0~95_combout  & ((\Mux29~11_combout  & ((\Mux3~8_combout ))) # (!\Mux29~11_combout  & (\Mux3~5_combout ))))

	.dataa(\Mux3~5_combout ),
	.datab(\Mux3~8_combout ),
	.datac(\Add0~95_combout ),
	.datad(\Mux29~11_combout ),
	.cin(gnd),
	.combout(Mux32),
	.cout());
// synopsys translate_off
defparam \Mux3~9 .lut_mask = 16'hCCCA;
defparam \Mux3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N24
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// Mux01 = (Mux0 & ((temp_ALUop_output_0) # (alu_a_mux_output_311))) # (!Mux0 & (temp_ALUop_output_0 & alu_a_mux_output_311))

	.dataa(Mux0),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(alu_a_mux_output_311),
	.cin(gnd),
	.combout(Mux01),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hFAA0;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N12
cycloneive_lcell_comb \Mux0~7 (
// Equation(s):
// Mux02 = (\Mux0~6_combout  & ((\Add0~103_combout ) # ((!\Mux19~1_combout )))) # (!\Mux0~6_combout  & (((\Mux0~5_combout  & \Mux19~1_combout ))))

	.dataa(\Add0~103_combout ),
	.datab(\Mux0~5_combout ),
	.datac(\Mux0~6_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(Mux02),
	.cout());
// synopsys translate_off
defparam \Mux0~7 .lut_mask = 16'hACF0;
defparam \Mux0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N26
cycloneive_lcell_comb \Mux1~2 (
// Equation(s):
// Mux110 = (alu_a_mux_output_30 & ((temp_ALUop_output_0) # (Mux1))) # (!alu_a_mux_output_30 & (temp_ALUop_output_0 & Mux1))

	.dataa(alu_a_mux_output_30),
	.datab(temp_ALUop_output_0),
	.datac(gnd),
	.datad(Mux1),
	.cin(gnd),
	.combout(Mux110),
	.cout());
// synopsys translate_off
defparam \Mux1~2 .lut_mask = 16'hEE88;
defparam \Mux1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N28
cycloneive_lcell_comb \Equal0~22 (
// Equation(s):
// Equal0 = (!Mux312 & (\Equal0~6_combout  & (\Equal0~10_combout  & \Equal0~21_combout )))

	.dataa(Mux312),
	.datab(\Equal0~6_combout ),
	.datac(\Equal0~10_combout ),
	.datad(\Equal0~21_combout ),
	.cin(gnd),
	.combout(Equal0),
	.cout());
// synopsys translate_off
defparam \Equal0~22 .lut_mask = 16'h4000;
defparam \Equal0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N18
cycloneive_lcell_comb \Mux1~10 (
// Equation(s):
// Mux113 = (\Mux1~9_combout  & ((\Mux1~7_combout ) # ((!\Mux19~1_combout )))) # (!\Mux1~9_combout  & (((\Add0~101_combout  & \Mux19~1_combout ))))

	.dataa(\Mux1~7_combout ),
	.datab(\Mux1~9_combout ),
	.datac(\Add0~101_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(Mux113),
	.cout());
// synopsys translate_off
defparam \Mux1~10 .lut_mask = 16'hB8CC;
defparam \Mux1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N18
cycloneive_lcell_comb \Mux5~8 (
// Equation(s):
// Mux51 = (\Mux5~7_combout  & ((\Mux5~5_combout ) # ((!\Mux19~1_combout )))) # (!\Mux5~7_combout  & (((\Mux19~1_combout  & \Add0~88_combout ))))

	.dataa(\Mux5~7_combout ),
	.datab(\Mux5~5_combout ),
	.datac(\Mux19~1_combout ),
	.datad(\Add0~88_combout ),
	.cin(gnd),
	.combout(Mux51),
	.cout());
// synopsys translate_off
defparam \Mux5~8 .lut_mask = 16'hDA8A;
defparam \Mux5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N6
cycloneive_lcell_comb \Mux7~7 (
// Equation(s):
// Mux71 = (\Mux7~6_combout  & ((\Mux7~5_combout ) # ((!\Mux19~1_combout )))) # (!\Mux7~6_combout  & (((\Mux19~1_combout  & \Add0~83_combout ))))

	.dataa(\Mux7~5_combout ),
	.datab(\Mux7~6_combout ),
	.datac(\Mux19~1_combout ),
	.datad(\Add0~83_combout ),
	.cin(gnd),
	.combout(Mux71),
	.cout());
// synopsys translate_off
defparam \Mux7~7 .lut_mask = 16'hBC8C;
defparam \Mux7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N0
cycloneive_lcell_comb \ShiftLeft0~13 (
// Equation(s):
// \ShiftLeft0~13_combout  = (Mux301) # ((Mux29) # ((!Mux16 & alu_b_mux_output_2)))

	.dataa(Mux301),
	.datab(Mux16),
	.datac(Mux29),
	.datad(alu_b_mux_output_2),
	.cin(gnd),
	.combout(\ShiftLeft0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~13 .lut_mask = 16'hFBFA;
defparam \ShiftLeft0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N22
cycloneive_lcell_comb \ShiftLeft0~12 (
// Equation(s):
// \ShiftLeft0~12_combout  = (Mux311 & ((alu_a_mux_output_0))) # (!Mux311 & (alu_a_mux_output_1))

	.dataa(alu_a_mux_output_1),
	.datab(gnd),
	.datac(alu_a_mux_output_0),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftLeft0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~12 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N0
cycloneive_lcell_comb \ShiftLeft0~14 (
// Equation(s):
// \ShiftLeft0~14_combout  = (!\ShiftLeft0~11_combout  & (!Mux281 & (!\ShiftLeft0~13_combout  & \ShiftLeft0~12_combout )))

	.dataa(\ShiftLeft0~11_combout ),
	.datab(Mux281),
	.datac(\ShiftLeft0~13_combout ),
	.datad(\ShiftLeft0~12_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~14 .lut_mask = 16'h0100;
defparam \ShiftLeft0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N20
cycloneive_lcell_comb \ShiftLeft0~15 (
// Equation(s):
// \ShiftLeft0~15_combout  = (!Mux271 & \ShiftLeft0~14_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux271),
	.datad(\ShiftLeft0~14_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~15 .lut_mask = 16'h0F00;
defparam \ShiftLeft0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N12
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (temp_ALUop_output_1 & (((temp_ALUop_output_0)))) # (!temp_ALUop_output_1 & ((temp_ALUop_output_0 & (\ShiftRight0~29_combout )) # (!temp_ALUop_output_0 & ((\ShiftLeft0~15_combout )))))

	.dataa(\ShiftRight0~29_combout ),
	.datab(temp_ALUop_output_1),
	.datac(temp_ALUop_output_0),
	.datad(\ShiftLeft0~15_combout ),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'hE3E0;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N6
cycloneive_lcell_comb \Mux30~3 (
// Equation(s):
// \Mux30~3_combout  = (\Mux30~2_combout  & (((alu_a_mux_output_1) # (Mux301)) # (!temp_ALUop_output_1))) # (!\Mux30~2_combout  & (temp_ALUop_output_1 & (alu_a_mux_output_1 & Mux301)))

	.dataa(\Mux30~2_combout ),
	.datab(temp_ALUop_output_1),
	.datac(alu_a_mux_output_1),
	.datad(Mux301),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~3 .lut_mask = 16'hEAA2;
defparam \Mux30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N18
cycloneive_lcell_comb \Add0~106 (
// Equation(s):
// \Add0~106_combout  = (!Mux31 & ((temp_ALUsrc_output_0 $ (temp_ALUsrc_output_1)) # (!alu_b_mux_output_01)))

	.dataa(Mux31),
	.datab(temp_ALUsrc_output_0),
	.datac(temp_ALUsrc_output_1),
	.datad(alu_b_mux_output_01),
	.cin(gnd),
	.combout(\Add0~106_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~106 .lut_mask = 16'h1455;
defparam \Add0~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N28
cycloneive_lcell_comb \Add0~5 (
// Equation(s):
// \Add0~5_combout  = temp_ALUop_output_0 $ ((((alu_b_mux_output_0 & !Mux16)) # (!\Add0~106_combout )))

	.dataa(temp_ALUop_output_0),
	.datab(\Add0~106_combout ),
	.datac(alu_b_mux_output_0),
	.datad(Mux16),
	.cin(gnd),
	.combout(\Add0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~5 .lut_mask = 16'h9959;
defparam \Add0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N16
cycloneive_lcell_comb \Add0~7 (
// Equation(s):
// \Add0~7_cout  = CARRY(temp_ALUop_output_0)

	.dataa(temp_ALUop_output_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add0~7_cout ));
// synopsys translate_off
defparam \Add0~7 .lut_mask = 16'h00AA;
defparam \Add0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N20
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = ((\Add0~4_combout  $ (alu_a_mux_output_1 $ (!\Add0~9 )))) # (GND)
// \Add0~11  = CARRY((\Add0~4_combout  & ((alu_a_mux_output_1) # (!\Add0~9 ))) # (!\Add0~4_combout  & (alu_a_mux_output_1 & !\Add0~9 )))

	.dataa(\Add0~4_combout ),
	.datab(alu_a_mux_output_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h698E;
defparam \Add0~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N28
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (!temp_ALUop_output_1 & ((temp_ALUop_output_0 & (!alu_a_mux_output_1 & !Mux301)) # (!temp_ALUop_output_0 & (alu_a_mux_output_1 $ (Mux301)))))

	.dataa(temp_ALUop_output_0),
	.datab(temp_ALUop_output_1),
	.datac(alu_a_mux_output_1),
	.datad(Mux301),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'h0112;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N18
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (\Mux30~0_combout ) # ((\Add0~10_combout  & temp_ALUop_output_1))

	.dataa(\Add0~10_combout ),
	.datab(temp_ALUop_output_1),
	.datac(gnd),
	.datad(\Mux30~0_combout ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hFF88;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N0
cycloneive_lcell_comb \LessThan0~1 (
// Equation(s):
// \LessThan0~1_cout  = CARRY((Mux311 & !alu_a_mux_output_0))

	.dataa(Mux311),
	.datab(alu_a_mux_output_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
// synopsys translate_off
defparam \LessThan0~1 .lut_mask = 16'h0022;
defparam \LessThan0~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N2
cycloneive_lcell_comb \LessThan0~3 (
// Equation(s):
// \LessThan0~3_cout  = CARRY((alu_a_mux_output_1 & ((!\LessThan0~1_cout ) # (!Mux301))) # (!alu_a_mux_output_1 & (!Mux301 & !\LessThan0~1_cout )))

	.dataa(alu_a_mux_output_1),
	.datab(Mux301),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
// synopsys translate_off
defparam \LessThan0~3 .lut_mask = 16'h002B;
defparam \LessThan0~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N4
cycloneive_lcell_comb \LessThan0~5 (
// Equation(s):
// \LessThan0~5_cout  = CARRY((alu_a_mux_output_2 & (Mux291 & !\LessThan0~3_cout )) # (!alu_a_mux_output_2 & ((Mux291) # (!\LessThan0~3_cout ))))

	.dataa(alu_a_mux_output_2),
	.datab(Mux291),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
// synopsys translate_off
defparam \LessThan0~5 .lut_mask = 16'h004D;
defparam \LessThan0~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N6
cycloneive_lcell_comb \LessThan0~7 (
// Equation(s):
// \LessThan0~7_cout  = CARRY((alu_a_mux_output_31 & ((!\LessThan0~5_cout ) # (!Mux281))) # (!alu_a_mux_output_31 & (!Mux281 & !\LessThan0~5_cout )))

	.dataa(alu_a_mux_output_31),
	.datab(Mux281),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
// synopsys translate_off
defparam \LessThan0~7 .lut_mask = 16'h002B;
defparam \LessThan0~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N8
cycloneive_lcell_comb \LessThan0~9 (
// Equation(s):
// \LessThan0~9_cout  = CARRY((Mux271 & ((!\LessThan0~7_cout ) # (!alu_a_mux_output_4))) # (!Mux271 & (!alu_a_mux_output_4 & !\LessThan0~7_cout )))

	.dataa(Mux271),
	.datab(alu_a_mux_output_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
// synopsys translate_off
defparam \LessThan0~9 .lut_mask = 16'h002B;
defparam \LessThan0~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N10
cycloneive_lcell_comb \LessThan0~11 (
// Equation(s):
// \LessThan0~11_cout  = CARRY((Mux26 & (alu_a_mux_output_5 & !\LessThan0~9_cout )) # (!Mux26 & ((alu_a_mux_output_5) # (!\LessThan0~9_cout ))))

	.dataa(Mux26),
	.datab(alu_a_mux_output_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
// synopsys translate_off
defparam \LessThan0~11 .lut_mask = 16'h004D;
defparam \LessThan0~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N12
cycloneive_lcell_comb \LessThan0~13 (
// Equation(s):
// \LessThan0~13_cout  = CARRY((Mux25 & ((!\LessThan0~11_cout ) # (!alu_a_mux_output_6))) # (!Mux25 & (!alu_a_mux_output_6 & !\LessThan0~11_cout )))

	.dataa(Mux25),
	.datab(alu_a_mux_output_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
// synopsys translate_off
defparam \LessThan0~13 .lut_mask = 16'h002B;
defparam \LessThan0~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N14
cycloneive_lcell_comb \LessThan0~15 (
// Equation(s):
// \LessThan0~15_cout  = CARRY((alu_a_mux_output_7 & ((!\LessThan0~13_cout ) # (!Mux24))) # (!alu_a_mux_output_7 & (!Mux24 & !\LessThan0~13_cout )))

	.dataa(alu_a_mux_output_7),
	.datab(Mux24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
// synopsys translate_off
defparam \LessThan0~15 .lut_mask = 16'h002B;
defparam \LessThan0~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N16
cycloneive_lcell_comb \LessThan0~17 (
// Equation(s):
// \LessThan0~17_cout  = CARRY((Mux23 & ((!\LessThan0~15_cout ) # (!alu_a_mux_output_8))) # (!Mux23 & (!alu_a_mux_output_8 & !\LessThan0~15_cout )))

	.dataa(Mux23),
	.datab(alu_a_mux_output_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~15_cout ),
	.combout(),
	.cout(\LessThan0~17_cout ));
// synopsys translate_off
defparam \LessThan0~17 .lut_mask = 16'h002B;
defparam \LessThan0~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N18
cycloneive_lcell_comb \LessThan0~19 (
// Equation(s):
// \LessThan0~19_cout  = CARRY((Mux22 & (alu_a_mux_output_9 & !\LessThan0~17_cout )) # (!Mux22 & ((alu_a_mux_output_9) # (!\LessThan0~17_cout ))))

	.dataa(Mux22),
	.datab(alu_a_mux_output_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~17_cout ),
	.combout(),
	.cout(\LessThan0~19_cout ));
// synopsys translate_off
defparam \LessThan0~19 .lut_mask = 16'h004D;
defparam \LessThan0~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N20
cycloneive_lcell_comb \LessThan0~21 (
// Equation(s):
// \LessThan0~21_cout  = CARRY((alu_a_mux_output_10 & (Mux21 & !\LessThan0~19_cout )) # (!alu_a_mux_output_10 & ((Mux21) # (!\LessThan0~19_cout ))))

	.dataa(alu_a_mux_output_10),
	.datab(Mux21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~19_cout ),
	.combout(),
	.cout(\LessThan0~21_cout ));
// synopsys translate_off
defparam \LessThan0~21 .lut_mask = 16'h004D;
defparam \LessThan0~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N22
cycloneive_lcell_comb \LessThan0~23 (
// Equation(s):
// \LessThan0~23_cout  = CARRY((Mux20 & (alu_a_mux_output_11 & !\LessThan0~21_cout )) # (!Mux20 & ((alu_a_mux_output_11) # (!\LessThan0~21_cout ))))

	.dataa(Mux20),
	.datab(alu_a_mux_output_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~21_cout ),
	.combout(),
	.cout(\LessThan0~23_cout ));
// synopsys translate_off
defparam \LessThan0~23 .lut_mask = 16'h004D;
defparam \LessThan0~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N24
cycloneive_lcell_comb \LessThan0~25 (
// Equation(s):
// \LessThan0~25_cout  = CARRY((Mux19 & ((!\LessThan0~23_cout ) # (!alu_a_mux_output_12))) # (!Mux19 & (!alu_a_mux_output_12 & !\LessThan0~23_cout )))

	.dataa(Mux19),
	.datab(alu_a_mux_output_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~23_cout ),
	.combout(),
	.cout(\LessThan0~25_cout ));
// synopsys translate_off
defparam \LessThan0~25 .lut_mask = 16'h002B;
defparam \LessThan0~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N26
cycloneive_lcell_comb \LessThan0~27 (
// Equation(s):
// \LessThan0~27_cout  = CARRY((Mux18 & (alu_a_mux_output_13 & !\LessThan0~25_cout )) # (!Mux18 & ((alu_a_mux_output_13) # (!\LessThan0~25_cout ))))

	.dataa(Mux18),
	.datab(alu_a_mux_output_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~25_cout ),
	.combout(),
	.cout(\LessThan0~27_cout ));
// synopsys translate_off
defparam \LessThan0~27 .lut_mask = 16'h004D;
defparam \LessThan0~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N28
cycloneive_lcell_comb \LessThan0~29 (
// Equation(s):
// \LessThan0~29_cout  = CARRY((Mux171 & ((!\LessThan0~27_cout ) # (!alu_a_mux_output_14))) # (!Mux171 & (!alu_a_mux_output_14 & !\LessThan0~27_cout )))

	.dataa(Mux171),
	.datab(alu_a_mux_output_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~27_cout ),
	.combout(),
	.cout(\LessThan0~29_cout ));
// synopsys translate_off
defparam \LessThan0~29 .lut_mask = 16'h002B;
defparam \LessThan0~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N30
cycloneive_lcell_comb \LessThan0~31 (
// Equation(s):
// \LessThan0~31_cout  = CARRY((Mux161 & (alu_a_mux_output_15 & !\LessThan0~29_cout )) # (!Mux161 & ((alu_a_mux_output_15) # (!\LessThan0~29_cout ))))

	.dataa(Mux161),
	.datab(alu_a_mux_output_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~29_cout ),
	.combout(),
	.cout(\LessThan0~31_cout ));
// synopsys translate_off
defparam \LessThan0~31 .lut_mask = 16'h004D;
defparam \LessThan0~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N0
cycloneive_lcell_comb \LessThan0~33 (
// Equation(s):
// \LessThan0~33_cout  = CARRY((alu_a_mux_output_16 & (Mux15 & !\LessThan0~31_cout )) # (!alu_a_mux_output_16 & ((Mux15) # (!\LessThan0~31_cout ))))

	.dataa(alu_a_mux_output_16),
	.datab(Mux15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~31_cout ),
	.combout(),
	.cout(\LessThan0~33_cout ));
// synopsys translate_off
defparam \LessThan0~33 .lut_mask = 16'h004D;
defparam \LessThan0~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N2
cycloneive_lcell_comb \LessThan0~35 (
// Equation(s):
// \LessThan0~35_cout  = CARRY((alu_a_mux_output_17 & ((!\LessThan0~33_cout ) # (!Mux14))) # (!alu_a_mux_output_17 & (!Mux14 & !\LessThan0~33_cout )))

	.dataa(alu_a_mux_output_17),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~33_cout ),
	.combout(),
	.cout(\LessThan0~35_cout ));
// synopsys translate_off
defparam \LessThan0~35 .lut_mask = 16'h002B;
defparam \LessThan0~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N4
cycloneive_lcell_comb \LessThan0~37 (
// Equation(s):
// \LessThan0~37_cout  = CARRY((alu_a_mux_output_18 & (Mux13 & !\LessThan0~35_cout )) # (!alu_a_mux_output_18 & ((Mux13) # (!\LessThan0~35_cout ))))

	.dataa(alu_a_mux_output_18),
	.datab(Mux13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~35_cout ),
	.combout(),
	.cout(\LessThan0~37_cout ));
// synopsys translate_off
defparam \LessThan0~37 .lut_mask = 16'h004D;
defparam \LessThan0~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N6
cycloneive_lcell_comb \LessThan0~39 (
// Equation(s):
// \LessThan0~39_cout  = CARRY((alu_a_mux_output_19 & ((!\LessThan0~37_cout ) # (!Mux12))) # (!alu_a_mux_output_19 & (!Mux12 & !\LessThan0~37_cout )))

	.dataa(alu_a_mux_output_19),
	.datab(Mux12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~37_cout ),
	.combout(),
	.cout(\LessThan0~39_cout ));
// synopsys translate_off
defparam \LessThan0~39 .lut_mask = 16'h002B;
defparam \LessThan0~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N8
cycloneive_lcell_comb \LessThan0~41 (
// Equation(s):
// \LessThan0~41_cout  = CARRY((Mux11 & ((!\LessThan0~39_cout ) # (!alu_a_mux_output_20))) # (!Mux11 & (!alu_a_mux_output_20 & !\LessThan0~39_cout )))

	.dataa(Mux11),
	.datab(alu_a_mux_output_20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~39_cout ),
	.combout(),
	.cout(\LessThan0~41_cout ));
// synopsys translate_off
defparam \LessThan0~41 .lut_mask = 16'h002B;
defparam \LessThan0~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N10
cycloneive_lcell_comb \LessThan0~43 (
// Equation(s):
// \LessThan0~43_cout  = CARRY((Mux10 & (alu_a_mux_output_21 & !\LessThan0~41_cout )) # (!Mux10 & ((alu_a_mux_output_21) # (!\LessThan0~41_cout ))))

	.dataa(Mux10),
	.datab(alu_a_mux_output_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~41_cout ),
	.combout(),
	.cout(\LessThan0~43_cout ));
// synopsys translate_off
defparam \LessThan0~43 .lut_mask = 16'h004D;
defparam \LessThan0~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N12
cycloneive_lcell_comb \LessThan0~45 (
// Equation(s):
// \LessThan0~45_cout  = CARRY((Mux9 & ((!\LessThan0~43_cout ) # (!alu_a_mux_output_22))) # (!Mux9 & (!alu_a_mux_output_22 & !\LessThan0~43_cout )))

	.dataa(Mux9),
	.datab(alu_a_mux_output_22),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~43_cout ),
	.combout(),
	.cout(\LessThan0~45_cout ));
// synopsys translate_off
defparam \LessThan0~45 .lut_mask = 16'h002B;
defparam \LessThan0~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N14
cycloneive_lcell_comb \LessThan0~47 (
// Equation(s):
// \LessThan0~47_cout  = CARRY((alu_a_mux_output_23 & ((!\LessThan0~45_cout ) # (!Mux8))) # (!alu_a_mux_output_23 & (!Mux8 & !\LessThan0~45_cout )))

	.dataa(alu_a_mux_output_23),
	.datab(Mux8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~45_cout ),
	.combout(),
	.cout(\LessThan0~47_cout ));
// synopsys translate_off
defparam \LessThan0~47 .lut_mask = 16'h002B;
defparam \LessThan0~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N16
cycloneive_lcell_comb \LessThan0~49 (
// Equation(s):
// \LessThan0~49_cout  = CARRY((alu_a_mux_output_24 & (Mux7 & !\LessThan0~47_cout )) # (!alu_a_mux_output_24 & ((Mux7) # (!\LessThan0~47_cout ))))

	.dataa(alu_a_mux_output_24),
	.datab(Mux7),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~47_cout ),
	.combout(),
	.cout(\LessThan0~49_cout ));
// synopsys translate_off
defparam \LessThan0~49 .lut_mask = 16'h004D;
defparam \LessThan0~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N18
cycloneive_lcell_comb \LessThan0~51 (
// Equation(s):
// \LessThan0~51_cout  = CARRY((Mux6 & (alu_a_mux_output_25 & !\LessThan0~49_cout )) # (!Mux6 & ((alu_a_mux_output_25) # (!\LessThan0~49_cout ))))

	.dataa(Mux6),
	.datab(alu_a_mux_output_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~49_cout ),
	.combout(),
	.cout(\LessThan0~51_cout ));
// synopsys translate_off
defparam \LessThan0~51 .lut_mask = 16'h004D;
defparam \LessThan0~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N20
cycloneive_lcell_comb \LessThan0~53 (
// Equation(s):
// \LessThan0~53_cout  = CARRY((Mux5 & ((!\LessThan0~51_cout ) # (!alu_a_mux_output_26))) # (!Mux5 & (!alu_a_mux_output_26 & !\LessThan0~51_cout )))

	.dataa(Mux5),
	.datab(alu_a_mux_output_26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~51_cout ),
	.combout(),
	.cout(\LessThan0~53_cout ));
// synopsys translate_off
defparam \LessThan0~53 .lut_mask = 16'h002B;
defparam \LessThan0~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N22
cycloneive_lcell_comb \LessThan0~55 (
// Equation(s):
// \LessThan0~55_cout  = CARRY((alu_a_mux_output_27 & ((!\LessThan0~53_cout ) # (!Mux4))) # (!alu_a_mux_output_27 & (!Mux4 & !\LessThan0~53_cout )))

	.dataa(alu_a_mux_output_27),
	.datab(Mux4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~53_cout ),
	.combout(),
	.cout(\LessThan0~55_cout ));
// synopsys translate_off
defparam \LessThan0~55 .lut_mask = 16'h002B;
defparam \LessThan0~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N24
cycloneive_lcell_comb \LessThan0~57 (
// Equation(s):
// \LessThan0~57_cout  = CARRY((alu_a_mux_output_28 & (Mux3 & !\LessThan0~55_cout )) # (!alu_a_mux_output_28 & ((Mux3) # (!\LessThan0~55_cout ))))

	.dataa(alu_a_mux_output_28),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~55_cout ),
	.combout(),
	.cout(\LessThan0~57_cout ));
// synopsys translate_off
defparam \LessThan0~57 .lut_mask = 16'h004D;
defparam \LessThan0~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N26
cycloneive_lcell_comb \LessThan0~59 (
// Equation(s):
// \LessThan0~59_cout  = CARRY((alu_a_mux_output_29 & ((!\LessThan0~57_cout ) # (!Mux2))) # (!alu_a_mux_output_29 & (!Mux2 & !\LessThan0~57_cout )))

	.dataa(alu_a_mux_output_29),
	.datab(Mux2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~57_cout ),
	.combout(),
	.cout(\LessThan0~59_cout ));
// synopsys translate_off
defparam \LessThan0~59 .lut_mask = 16'h002B;
defparam \LessThan0~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N28
cycloneive_lcell_comb \LessThan0~61 (
// Equation(s):
// \LessThan0~61_cout  = CARRY((alu_a_mux_output_30 & (Mux1 & !\LessThan0~59_cout )) # (!alu_a_mux_output_30 & ((Mux1) # (!\LessThan0~59_cout ))))

	.dataa(alu_a_mux_output_30),
	.datab(Mux1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~59_cout ),
	.combout(),
	.cout(\LessThan0~61_cout ));
// synopsys translate_off
defparam \LessThan0~61 .lut_mask = 16'h004D;
defparam \LessThan0~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N30
cycloneive_lcell_comb \LessThan0~62 (
// Equation(s):
// \LessThan0~62_combout  = (Mux0 & (\LessThan0~61_cout  & alu_a_mux_output_311)) # (!Mux0 & ((\LessThan0~61_cout ) # (alu_a_mux_output_311)))

	.dataa(gnd),
	.datab(Mux0),
	.datac(gnd),
	.datad(alu_a_mux_output_311),
	.cin(\LessThan0~61_cout ),
	.combout(\LessThan0~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan0~62 .lut_mask = 16'hF330;
defparam \LessThan0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N0
cycloneive_lcell_comb \LessThan1~1 (
// Equation(s):
// \LessThan1~1_cout  = CARRY((Mux311 & !alu_a_mux_output_0))

	.dataa(Mux311),
	.datab(alu_a_mux_output_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan1~1_cout ));
// synopsys translate_off
defparam \LessThan1~1 .lut_mask = 16'h0022;
defparam \LessThan1~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N2
cycloneive_lcell_comb \LessThan1~3 (
// Equation(s):
// \LessThan1~3_cout  = CARRY((Mux301 & (alu_a_mux_output_1 & !\LessThan1~1_cout )) # (!Mux301 & ((alu_a_mux_output_1) # (!\LessThan1~1_cout ))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~1_cout ),
	.combout(),
	.cout(\LessThan1~3_cout ));
// synopsys translate_off
defparam \LessThan1~3 .lut_mask = 16'h004D;
defparam \LessThan1~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N4
cycloneive_lcell_comb \LessThan1~5 (
// Equation(s):
// \LessThan1~5_cout  = CARRY((alu_a_mux_output_2 & (Mux291 & !\LessThan1~3_cout )) # (!alu_a_mux_output_2 & ((Mux291) # (!\LessThan1~3_cout ))))

	.dataa(alu_a_mux_output_2),
	.datab(Mux291),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~3_cout ),
	.combout(),
	.cout(\LessThan1~5_cout ));
// synopsys translate_off
defparam \LessThan1~5 .lut_mask = 16'h004D;
defparam \LessThan1~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N6
cycloneive_lcell_comb \LessThan1~7 (
// Equation(s):
// \LessThan1~7_cout  = CARRY((Mux281 & (alu_a_mux_output_31 & !\LessThan1~5_cout )) # (!Mux281 & ((alu_a_mux_output_31) # (!\LessThan1~5_cout ))))

	.dataa(Mux281),
	.datab(alu_a_mux_output_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~5_cout ),
	.combout(),
	.cout(\LessThan1~7_cout ));
// synopsys translate_off
defparam \LessThan1~7 .lut_mask = 16'h004D;
defparam \LessThan1~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N8
cycloneive_lcell_comb \LessThan1~9 (
// Equation(s):
// \LessThan1~9_cout  = CARRY((Mux271 & ((!\LessThan1~7_cout ) # (!alu_a_mux_output_4))) # (!Mux271 & (!alu_a_mux_output_4 & !\LessThan1~7_cout )))

	.dataa(Mux271),
	.datab(alu_a_mux_output_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~7_cout ),
	.combout(),
	.cout(\LessThan1~9_cout ));
// synopsys translate_off
defparam \LessThan1~9 .lut_mask = 16'h002B;
defparam \LessThan1~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N10
cycloneive_lcell_comb \LessThan1~11 (
// Equation(s):
// \LessThan1~11_cout  = CARRY((Mux26 & (alu_a_mux_output_5 & !\LessThan1~9_cout )) # (!Mux26 & ((alu_a_mux_output_5) # (!\LessThan1~9_cout ))))

	.dataa(Mux26),
	.datab(alu_a_mux_output_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~9_cout ),
	.combout(),
	.cout(\LessThan1~11_cout ));
// synopsys translate_off
defparam \LessThan1~11 .lut_mask = 16'h004D;
defparam \LessThan1~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N12
cycloneive_lcell_comb \LessThan1~13 (
// Equation(s):
// \LessThan1~13_cout  = CARRY((Mux25 & ((!\LessThan1~11_cout ) # (!alu_a_mux_output_6))) # (!Mux25 & (!alu_a_mux_output_6 & !\LessThan1~11_cout )))

	.dataa(Mux25),
	.datab(alu_a_mux_output_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~11_cout ),
	.combout(),
	.cout(\LessThan1~13_cout ));
// synopsys translate_off
defparam \LessThan1~13 .lut_mask = 16'h002B;
defparam \LessThan1~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N14
cycloneive_lcell_comb \LessThan1~15 (
// Equation(s):
// \LessThan1~15_cout  = CARRY((Mux24 & (alu_a_mux_output_7 & !\LessThan1~13_cout )) # (!Mux24 & ((alu_a_mux_output_7) # (!\LessThan1~13_cout ))))

	.dataa(Mux24),
	.datab(alu_a_mux_output_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~13_cout ),
	.combout(),
	.cout(\LessThan1~15_cout ));
// synopsys translate_off
defparam \LessThan1~15 .lut_mask = 16'h004D;
defparam \LessThan1~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N16
cycloneive_lcell_comb \LessThan1~17 (
// Equation(s):
// \LessThan1~17_cout  = CARRY((Mux23 & ((!\LessThan1~15_cout ) # (!alu_a_mux_output_8))) # (!Mux23 & (!alu_a_mux_output_8 & !\LessThan1~15_cout )))

	.dataa(Mux23),
	.datab(alu_a_mux_output_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~15_cout ),
	.combout(),
	.cout(\LessThan1~17_cout ));
// synopsys translate_off
defparam \LessThan1~17 .lut_mask = 16'h002B;
defparam \LessThan1~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N18
cycloneive_lcell_comb \LessThan1~19 (
// Equation(s):
// \LessThan1~19_cout  = CARRY((alu_a_mux_output_9 & ((!\LessThan1~17_cout ) # (!Mux22))) # (!alu_a_mux_output_9 & (!Mux22 & !\LessThan1~17_cout )))

	.dataa(alu_a_mux_output_9),
	.datab(Mux22),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~17_cout ),
	.combout(),
	.cout(\LessThan1~19_cout ));
// synopsys translate_off
defparam \LessThan1~19 .lut_mask = 16'h002B;
defparam \LessThan1~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N20
cycloneive_lcell_comb \LessThan1~21 (
// Equation(s):
// \LessThan1~21_cout  = CARRY((Mux21 & ((!\LessThan1~19_cout ) # (!alu_a_mux_output_10))) # (!Mux21 & (!alu_a_mux_output_10 & !\LessThan1~19_cout )))

	.dataa(Mux21),
	.datab(alu_a_mux_output_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~19_cout ),
	.combout(),
	.cout(\LessThan1~21_cout ));
// synopsys translate_off
defparam \LessThan1~21 .lut_mask = 16'h002B;
defparam \LessThan1~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N22
cycloneive_lcell_comb \LessThan1~23 (
// Equation(s):
// \LessThan1~23_cout  = CARRY((alu_a_mux_output_11 & ((!\LessThan1~21_cout ) # (!Mux20))) # (!alu_a_mux_output_11 & (!Mux20 & !\LessThan1~21_cout )))

	.dataa(alu_a_mux_output_11),
	.datab(Mux20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~21_cout ),
	.combout(),
	.cout(\LessThan1~23_cout ));
// synopsys translate_off
defparam \LessThan1~23 .lut_mask = 16'h002B;
defparam \LessThan1~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N24
cycloneive_lcell_comb \LessThan1~25 (
// Equation(s):
// \LessThan1~25_cout  = CARRY((alu_a_mux_output_12 & (Mux19 & !\LessThan1~23_cout )) # (!alu_a_mux_output_12 & ((Mux19) # (!\LessThan1~23_cout ))))

	.dataa(alu_a_mux_output_12),
	.datab(Mux19),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~23_cout ),
	.combout(),
	.cout(\LessThan1~25_cout ));
// synopsys translate_off
defparam \LessThan1~25 .lut_mask = 16'h004D;
defparam \LessThan1~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N26
cycloneive_lcell_comb \LessThan1~27 (
// Equation(s):
// \LessThan1~27_cout  = CARRY((Mux18 & (alu_a_mux_output_13 & !\LessThan1~25_cout )) # (!Mux18 & ((alu_a_mux_output_13) # (!\LessThan1~25_cout ))))

	.dataa(Mux18),
	.datab(alu_a_mux_output_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~25_cout ),
	.combout(),
	.cout(\LessThan1~27_cout ));
// synopsys translate_off
defparam \LessThan1~27 .lut_mask = 16'h004D;
defparam \LessThan1~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N28
cycloneive_lcell_comb \LessThan1~29 (
// Equation(s):
// \LessThan1~29_cout  = CARRY((alu_a_mux_output_14 & (Mux171 & !\LessThan1~27_cout )) # (!alu_a_mux_output_14 & ((Mux171) # (!\LessThan1~27_cout ))))

	.dataa(alu_a_mux_output_14),
	.datab(Mux171),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~27_cout ),
	.combout(),
	.cout(\LessThan1~29_cout ));
// synopsys translate_off
defparam \LessThan1~29 .lut_mask = 16'h004D;
defparam \LessThan1~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N30
cycloneive_lcell_comb \LessThan1~31 (
// Equation(s):
// \LessThan1~31_cout  = CARRY((alu_a_mux_output_15 & ((!\LessThan1~29_cout ) # (!Mux161))) # (!alu_a_mux_output_15 & (!Mux161 & !\LessThan1~29_cout )))

	.dataa(alu_a_mux_output_15),
	.datab(Mux161),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~29_cout ),
	.combout(),
	.cout(\LessThan1~31_cout ));
// synopsys translate_off
defparam \LessThan1~31 .lut_mask = 16'h002B;
defparam \LessThan1~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N0
cycloneive_lcell_comb \LessThan1~33 (
// Equation(s):
// \LessThan1~33_cout  = CARRY((alu_a_mux_output_16 & (Mux15 & !\LessThan1~31_cout )) # (!alu_a_mux_output_16 & ((Mux15) # (!\LessThan1~31_cout ))))

	.dataa(alu_a_mux_output_16),
	.datab(Mux15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~31_cout ),
	.combout(),
	.cout(\LessThan1~33_cout ));
// synopsys translate_off
defparam \LessThan1~33 .lut_mask = 16'h004D;
defparam \LessThan1~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N2
cycloneive_lcell_comb \LessThan1~35 (
// Equation(s):
// \LessThan1~35_cout  = CARRY((Mux14 & (alu_a_mux_output_17 & !\LessThan1~33_cout )) # (!Mux14 & ((alu_a_mux_output_17) # (!\LessThan1~33_cout ))))

	.dataa(Mux14),
	.datab(alu_a_mux_output_17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~33_cout ),
	.combout(),
	.cout(\LessThan1~35_cout ));
// synopsys translate_off
defparam \LessThan1~35 .lut_mask = 16'h004D;
defparam \LessThan1~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N4
cycloneive_lcell_comb \LessThan1~37 (
// Equation(s):
// \LessThan1~37_cout  = CARRY((Mux13 & ((!\LessThan1~35_cout ) # (!alu_a_mux_output_18))) # (!Mux13 & (!alu_a_mux_output_18 & !\LessThan1~35_cout )))

	.dataa(Mux13),
	.datab(alu_a_mux_output_18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~35_cout ),
	.combout(),
	.cout(\LessThan1~37_cout ));
// synopsys translate_off
defparam \LessThan1~37 .lut_mask = 16'h002B;
defparam \LessThan1~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N6
cycloneive_lcell_comb \LessThan1~39 (
// Equation(s):
// \LessThan1~39_cout  = CARRY((Mux12 & (alu_a_mux_output_19 & !\LessThan1~37_cout )) # (!Mux12 & ((alu_a_mux_output_19) # (!\LessThan1~37_cout ))))

	.dataa(Mux12),
	.datab(alu_a_mux_output_19),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~37_cout ),
	.combout(),
	.cout(\LessThan1~39_cout ));
// synopsys translate_off
defparam \LessThan1~39 .lut_mask = 16'h004D;
defparam \LessThan1~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N8
cycloneive_lcell_comb \LessThan1~41 (
// Equation(s):
// \LessThan1~41_cout  = CARRY((alu_a_mux_output_20 & (Mux11 & !\LessThan1~39_cout )) # (!alu_a_mux_output_20 & ((Mux11) # (!\LessThan1~39_cout ))))

	.dataa(alu_a_mux_output_20),
	.datab(Mux11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~39_cout ),
	.combout(),
	.cout(\LessThan1~41_cout ));
// synopsys translate_off
defparam \LessThan1~41 .lut_mask = 16'h004D;
defparam \LessThan1~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N10
cycloneive_lcell_comb \LessThan1~43 (
// Equation(s):
// \LessThan1~43_cout  = CARRY((alu_a_mux_output_21 & ((!\LessThan1~41_cout ) # (!Mux10))) # (!alu_a_mux_output_21 & (!Mux10 & !\LessThan1~41_cout )))

	.dataa(alu_a_mux_output_21),
	.datab(Mux10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~41_cout ),
	.combout(),
	.cout(\LessThan1~43_cout ));
// synopsys translate_off
defparam \LessThan1~43 .lut_mask = 16'h002B;
defparam \LessThan1~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N12
cycloneive_lcell_comb \LessThan1~45 (
// Equation(s):
// \LessThan1~45_cout  = CARRY((alu_a_mux_output_22 & (Mux9 & !\LessThan1~43_cout )) # (!alu_a_mux_output_22 & ((Mux9) # (!\LessThan1~43_cout ))))

	.dataa(alu_a_mux_output_22),
	.datab(Mux9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~43_cout ),
	.combout(),
	.cout(\LessThan1~45_cout ));
// synopsys translate_off
defparam \LessThan1~45 .lut_mask = 16'h004D;
defparam \LessThan1~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N14
cycloneive_lcell_comb \LessThan1~47 (
// Equation(s):
// \LessThan1~47_cout  = CARRY((Mux8 & (alu_a_mux_output_23 & !\LessThan1~45_cout )) # (!Mux8 & ((alu_a_mux_output_23) # (!\LessThan1~45_cout ))))

	.dataa(Mux8),
	.datab(alu_a_mux_output_23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~45_cout ),
	.combout(),
	.cout(\LessThan1~47_cout ));
// synopsys translate_off
defparam \LessThan1~47 .lut_mask = 16'h004D;
defparam \LessThan1~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N16
cycloneive_lcell_comb \LessThan1~49 (
// Equation(s):
// \LessThan1~49_cout  = CARRY((Mux7 & ((!\LessThan1~47_cout ) # (!alu_a_mux_output_24))) # (!Mux7 & (!alu_a_mux_output_24 & !\LessThan1~47_cout )))

	.dataa(Mux7),
	.datab(alu_a_mux_output_24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~47_cout ),
	.combout(),
	.cout(\LessThan1~49_cout ));
// synopsys translate_off
defparam \LessThan1~49 .lut_mask = 16'h002B;
defparam \LessThan1~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N18
cycloneive_lcell_comb \LessThan1~51 (
// Equation(s):
// \LessThan1~51_cout  = CARRY((Mux6 & (alu_a_mux_output_25 & !\LessThan1~49_cout )) # (!Mux6 & ((alu_a_mux_output_25) # (!\LessThan1~49_cout ))))

	.dataa(Mux6),
	.datab(alu_a_mux_output_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~49_cout ),
	.combout(),
	.cout(\LessThan1~51_cout ));
// synopsys translate_off
defparam \LessThan1~51 .lut_mask = 16'h004D;
defparam \LessThan1~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N20
cycloneive_lcell_comb \LessThan1~53 (
// Equation(s):
// \LessThan1~53_cout  = CARRY((Mux5 & ((!\LessThan1~51_cout ) # (!alu_a_mux_output_26))) # (!Mux5 & (!alu_a_mux_output_26 & !\LessThan1~51_cout )))

	.dataa(Mux5),
	.datab(alu_a_mux_output_26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~51_cout ),
	.combout(),
	.cout(\LessThan1~53_cout ));
// synopsys translate_off
defparam \LessThan1~53 .lut_mask = 16'h002B;
defparam \LessThan1~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N22
cycloneive_lcell_comb \LessThan1~55 (
// Equation(s):
// \LessThan1~55_cout  = CARRY((Mux4 & (alu_a_mux_output_27 & !\LessThan1~53_cout )) # (!Mux4 & ((alu_a_mux_output_27) # (!\LessThan1~53_cout ))))

	.dataa(Mux4),
	.datab(alu_a_mux_output_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~53_cout ),
	.combout(),
	.cout(\LessThan1~55_cout ));
// synopsys translate_off
defparam \LessThan1~55 .lut_mask = 16'h004D;
defparam \LessThan1~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N24
cycloneive_lcell_comb \LessThan1~57 (
// Equation(s):
// \LessThan1~57_cout  = CARRY((alu_a_mux_output_28 & (Mux3 & !\LessThan1~55_cout )) # (!alu_a_mux_output_28 & ((Mux3) # (!\LessThan1~55_cout ))))

	.dataa(alu_a_mux_output_28),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~55_cout ),
	.combout(),
	.cout(\LessThan1~57_cout ));
// synopsys translate_off
defparam \LessThan1~57 .lut_mask = 16'h004D;
defparam \LessThan1~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N26
cycloneive_lcell_comb \LessThan1~59 (
// Equation(s):
// \LessThan1~59_cout  = CARRY((alu_a_mux_output_29 & ((!\LessThan1~57_cout ) # (!Mux2))) # (!alu_a_mux_output_29 & (!Mux2 & !\LessThan1~57_cout )))

	.dataa(alu_a_mux_output_29),
	.datab(Mux2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~57_cout ),
	.combout(),
	.cout(\LessThan1~59_cout ));
// synopsys translate_off
defparam \LessThan1~59 .lut_mask = 16'h002B;
defparam \LessThan1~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N28
cycloneive_lcell_comb \LessThan1~61 (
// Equation(s):
// \LessThan1~61_cout  = CARRY((alu_a_mux_output_30 & (Mux1 & !\LessThan1~59_cout )) # (!alu_a_mux_output_30 & ((Mux1) # (!\LessThan1~59_cout ))))

	.dataa(alu_a_mux_output_30),
	.datab(Mux1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~59_cout ),
	.combout(),
	.cout(\LessThan1~61_cout ));
// synopsys translate_off
defparam \LessThan1~61 .lut_mask = 16'h004D;
defparam \LessThan1~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N30
cycloneive_lcell_comb \LessThan1~62 (
// Equation(s):
// \LessThan1~62_combout  = (Mux0 & ((\LessThan1~61_cout ) # (!alu_a_mux_output_311))) # (!Mux0 & (\LessThan1~61_cout  & !alu_a_mux_output_311))

	.dataa(gnd),
	.datab(Mux0),
	.datac(gnd),
	.datad(alu_a_mux_output_311),
	.cin(\LessThan1~61_cout ),
	.combout(\LessThan1~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan1~62 .lut_mask = 16'hC0FC;
defparam \LessThan1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N6
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (temp_ALUop_output_0 & ((Mux311) # (alu_a_mux_output_0))) # (!temp_ALUop_output_0 & (Mux311 & alu_a_mux_output_0))

	.dataa(temp_ALUop_output_0),
	.datab(gnd),
	.datac(Mux311),
	.datad(alu_a_mux_output_0),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hFAA0;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N2
cycloneive_lcell_comb \Mux31~6 (
// Equation(s):
// \Mux31~6_combout  = (temp_ALUop_output_1 & (((\Mux31~2_combout ) # (temp_ALUop_output_3)))) # (!temp_ALUop_output_1 & (\Mux31~5_combout  & ((!temp_ALUop_output_3))))

	.dataa(\Mux31~5_combout ),
	.datab(temp_ALUop_output_1),
	.datac(\Mux31~2_combout ),
	.datad(temp_ALUop_output_3),
	.cin(gnd),
	.combout(\Mux31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~6 .lut_mask = 16'hCCE2;
defparam \Mux31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N24
cycloneive_lcell_comb \Mux31~7 (
// Equation(s):
// \Mux31~7_combout  = (temp_ALUop_output_2 & (\Mux31~1_combout  & ((!temp_ALUop_output_3)))) # (!temp_ALUop_output_2 & ((\Mux31~6_combout  $ (temp_ALUop_output_3))))

	.dataa(\Mux31~1_combout ),
	.datab(\Mux31~6_combout ),
	.datac(temp_ALUop_output_2),
	.datad(temp_ALUop_output_3),
	.cin(gnd),
	.combout(\Mux31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~7 .lut_mask = 16'h03AC;
defparam \Mux31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N6
cycloneive_lcell_comb \Mux31~8 (
// Equation(s):
// \Mux31~8_combout  = (\Mux31~7_combout  & ((\LessThan1~62_combout ) # ((!temp_ALUop_output_0) # (!temp_ALUop_output_3))))

	.dataa(\LessThan1~62_combout ),
	.datab(temp_ALUop_output_3),
	.datac(temp_ALUop_output_0),
	.datad(\Mux31~7_combout ),
	.cin(gnd),
	.combout(\Mux31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~8 .lut_mask = 16'hBF00;
defparam \Mux31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N2
cycloneive_lcell_comb \Mux29~11 (
// Equation(s):
// \Mux29~11_combout  = (!temp_ALUop_output_2 & (temp_ALUop_output_0 & temp_ALUop_output_1))

	.dataa(temp_ALUop_output_2),
	.datab(temp_ALUop_output_0),
	.datac(gnd),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Mux29~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~11 .lut_mask = 16'h4400;
defparam \Mux29~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N0
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (temp_ALUop_output_1) # (!temp_ALUop_output_2)

	.dataa(temp_ALUop_output_2),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hFF55;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N14
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (Mux281) # ((!Mux291 & Mux301))

	.dataa(gnd),
	.datab(Mux291),
	.datac(Mux301),
	.datad(Mux281),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hFF30;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N20
cycloneive_lcell_comb \ShiftRight0~34 (
// Equation(s):
// \ShiftRight0~34_combout  = (Mux311 & ((alu_a_mux_output_5))) # (!Mux311 & (alu_a_mux_output_4))

	.dataa(Mux311),
	.datab(gnd),
	.datac(alu_a_mux_output_4),
	.datad(alu_a_mux_output_5),
	.cin(gnd),
	.combout(\ShiftRight0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~34 .lut_mask = 16'hFA50;
defparam \ShiftRight0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N26
cycloneive_lcell_comb \ShiftRight0~57 (
// Equation(s):
// \ShiftRight0~57_combout  = (Mux301 & ((alu_a_mux_output_9))) # (!Mux301 & (alu_a_mux_output_7))

	.dataa(gnd),
	.datab(Mux301),
	.datac(alu_a_mux_output_7),
	.datad(alu_a_mux_output_9),
	.cin(gnd),
	.combout(\ShiftRight0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~57 .lut_mask = 16'hFC30;
defparam \ShiftRight0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N28
cycloneive_lcell_comb \ShiftRight0~56 (
// Equation(s):
// \ShiftRight0~56_combout  = (!Mux311 & ((Mux301 & (alu_a_mux_output_8)) # (!Mux301 & ((alu_a_mux_output_6)))))

	.dataa(alu_a_mux_output_8),
	.datab(Mux311),
	.datac(Mux301),
	.datad(alu_a_mux_output_6),
	.cin(gnd),
	.combout(\ShiftRight0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~56 .lut_mask = 16'h2320;
defparam \ShiftRight0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N8
cycloneive_lcell_comb \ShiftRight0~58 (
// Equation(s):
// \ShiftRight0~58_combout  = (\ShiftRight0~56_combout ) # ((Mux311 & \ShiftRight0~57_combout ))

	.dataa(Mux311),
	.datab(gnd),
	.datac(\ShiftRight0~57_combout ),
	.datad(\ShiftRight0~56_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~58 .lut_mask = 16'hFFA0;
defparam \ShiftRight0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N12
cycloneive_lcell_comb \ShiftRight0~31 (
// Equation(s):
// \ShiftRight0~31_combout  = (Mux311 & (alu_a_mux_output_31)) # (!Mux311 & ((alu_a_mux_output_2)))

	.dataa(gnd),
	.datab(Mux311),
	.datac(alu_a_mux_output_31),
	.datad(alu_a_mux_output_2),
	.cin(gnd),
	.combout(\ShiftRight0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~31 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N20
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (\ShiftRight0~59_combout  & (((!\Mux29~0_combout  & \ShiftRight0~31_combout )))) # (!\ShiftRight0~59_combout  & ((\ShiftRight0~58_combout ) # ((\Mux29~0_combout ))))

	.dataa(\ShiftRight0~59_combout ),
	.datab(\ShiftRight0~58_combout ),
	.datac(\Mux29~0_combout ),
	.datad(\ShiftRight0~31_combout ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'h5E54;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N24
cycloneive_lcell_comb \Mux29~2 (
// Equation(s):
// \Mux29~2_combout  = (\Mux29~0_combout  & ((\Mux29~1_combout  & (\ShiftRight0~64_combout )) # (!\Mux29~1_combout  & ((\ShiftRight0~34_combout ))))) # (!\Mux29~0_combout  & (((\Mux29~1_combout ))))

	.dataa(\ShiftRight0~64_combout ),
	.datab(\Mux29~0_combout ),
	.datac(\ShiftRight0~34_combout ),
	.datad(\Mux29~1_combout ),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~2 .lut_mask = 16'hBBC0;
defparam \Mux29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N26
cycloneive_lcell_comb \ShiftRight0~71 (
// Equation(s):
// \ShiftRight0~71_combout  = (Mux301 & ((Mux311 & (alu_a_mux_output_21)) # (!Mux311 & ((alu_a_mux_output_20)))))

	.dataa(alu_a_mux_output_21),
	.datab(Mux311),
	.datac(Mux301),
	.datad(alu_a_mux_output_20),
	.cin(gnd),
	.combout(\ShiftRight0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~71 .lut_mask = 16'hB080;
defparam \ShiftRight0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N8
cycloneive_lcell_comb \ShiftRight0~72 (
// Equation(s):
// \ShiftRight0~72_combout  = (!Mux301 & ((Mux311 & ((alu_a_mux_output_19))) # (!Mux311 & (alu_a_mux_output_18))))

	.dataa(alu_a_mux_output_18),
	.datab(Mux311),
	.datac(Mux301),
	.datad(alu_a_mux_output_19),
	.cin(gnd),
	.combout(\ShiftRight0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~72 .lut_mask = 16'h0E02;
defparam \ShiftRight0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N4
cycloneive_lcell_comb \ShiftRight0~73 (
// Equation(s):
// \ShiftRight0~73_combout  = (Mux291 & (\ShiftRight0~70_combout )) # (!Mux291 & (((\ShiftRight0~71_combout ) # (\ShiftRight0~72_combout ))))

	.dataa(\ShiftRight0~70_combout ),
	.datab(Mux291),
	.datac(\ShiftRight0~71_combout ),
	.datad(\ShiftRight0~72_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~73 .lut_mask = 16'hBBB8;
defparam \ShiftRight0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N4
cycloneive_lcell_comb \ShiftRight0~65 (
// Equation(s):
// \ShiftRight0~65_combout  = (Mux311 & ((Mux301 & (alu_a_mux_output_29)) # (!Mux301 & ((alu_a_mux_output_27)))))

	.dataa(Mux311),
	.datab(alu_a_mux_output_29),
	.datac(alu_a_mux_output_27),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftRight0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~65 .lut_mask = 16'h88A0;
defparam \ShiftRight0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N24
cycloneive_lcell_comb \ShiftRight0~66 (
// Equation(s):
// \ShiftRight0~66_combout  = (!Mux311 & ((Mux301 & (alu_a_mux_output_28)) # (!Mux301 & ((alu_a_mux_output_26)))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_28),
	.datac(Mux311),
	.datad(alu_a_mux_output_26),
	.cin(gnd),
	.combout(\ShiftRight0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~66 .lut_mask = 16'h0D08;
defparam \ShiftRight0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N18
cycloneive_lcell_comb \ShiftRight0~67 (
// Equation(s):
// \ShiftRight0~67_combout  = (!Mux291 & ((\ShiftRight0~65_combout ) # (\ShiftRight0~66_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~65_combout ),
	.datac(Mux291),
	.datad(\ShiftRight0~66_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~67 .lut_mask = 16'h0F0C;
defparam \ShiftRight0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N8
cycloneive_lcell_comb \ShiftRight0~44 (
// Equation(s):
// \ShiftRight0~44_combout  = (Mux311 & ((alu_a_mux_output_311))) # (!Mux311 & (alu_a_mux_output_30))

	.dataa(gnd),
	.datab(alu_a_mux_output_30),
	.datac(alu_a_mux_output_311),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftRight0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~44 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N24
cycloneive_lcell_comb \ShiftRight0~68 (
// Equation(s):
// \ShiftRight0~68_combout  = (\ShiftRight0~67_combout ) # ((!Mux301 & (Mux291 & \ShiftRight0~44_combout )))

	.dataa(Mux301),
	.datab(\ShiftRight0~67_combout ),
	.datac(Mux291),
	.datad(\ShiftRight0~44_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~68 .lut_mask = 16'hDCCC;
defparam \ShiftRight0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N14
cycloneive_lcell_comb \ShiftRight0~74 (
// Equation(s):
// \ShiftRight0~74_combout  = (Mux281 & ((\ShiftRight0~68_combout ))) # (!Mux281 & (\ShiftRight0~73_combout ))

	.dataa(Mux281),
	.datab(gnd),
	.datac(\ShiftRight0~73_combout ),
	.datad(\ShiftRight0~68_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~74 .lut_mask = 16'hFA50;
defparam \ShiftRight0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N8
cycloneive_lcell_comb \Mux29~3 (
// Equation(s):
// \Mux29~3_combout  = (temp_ALUop_output_0 & !temp_ALUop_output_1)

	.dataa(gnd),
	.datab(temp_ALUop_output_0),
	.datac(temp_ALUop_output_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~3 .lut_mask = 16'h0C0C;
defparam \Mux29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N30
cycloneive_lcell_comb \Mux29~7 (
// Equation(s):
// \Mux29~7_combout  = (\Mux29~6_combout  & (((\ShiftRight0~74_combout ) # (!\Mux29~3_combout )))) # (!\Mux29~6_combout  & (\Mux29~2_combout  & ((\Mux29~3_combout ))))

	.dataa(\Mux29~6_combout ),
	.datab(\Mux29~2_combout ),
	.datac(\ShiftRight0~74_combout ),
	.datad(\Mux29~3_combout ),
	.cin(gnd),
	.combout(\Mux29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~7 .lut_mask = 16'hE4AA;
defparam \Mux29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N10
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (temp_ALUop_output_2 & ((temp_ALUop_output_0) # (temp_ALUop_output_1)))

	.dataa(temp_ALUop_output_0),
	.datab(temp_ALUop_output_2),
	.datac(gnd),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hCC88;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N20
cycloneive_lcell_comb \ShiftLeft0~9 (
// Equation(s):
// \ShiftLeft0~9_combout  = (Mux23) # ((Mux25) # ((Mux22) # (Mux24)))

	.dataa(Mux23),
	.datab(Mux25),
	.datac(Mux22),
	.datad(Mux24),
	.cin(gnd),
	.combout(\ShiftLeft0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~9 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N14
cycloneive_lcell_comb \ShiftLeft0~10 (
// Equation(s):
// \ShiftLeft0~10_combout  = (Mux18) # ((Mux26) # ((Mux20) # (\ShiftLeft0~9_combout )))

	.dataa(Mux18),
	.datab(Mux26),
	.datac(Mux20),
	.datad(\ShiftLeft0~9_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~10 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N2
cycloneive_lcell_comb \ShiftLeft0~4 (
// Equation(s):
// \ShiftLeft0~4_combout  = (Mux5) # ((Mux6) # ((Mux8) # (Mux7)))

	.dataa(Mux5),
	.datab(Mux6),
	.datac(Mux8),
	.datad(Mux7),
	.cin(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~4 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N22
cycloneive_lcell_comb \ShiftLeft0~2 (
// Equation(s):
// \ShiftLeft0~2_combout  = (Mux13) # ((Mux14) # ((Mux15) # (Mux4)))

	.dataa(Mux13),
	.datab(Mux14),
	.datac(Mux15),
	.datad(Mux4),
	.cin(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~2 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N16
cycloneive_lcell_comb \ShiftLeft0~3 (
// Equation(s):
// \ShiftLeft0~3_combout  = (Mux3) # ((Mux0) # ((Mux2) # (Mux1)))

	.dataa(Mux3),
	.datab(Mux0),
	.datac(Mux2),
	.datad(Mux1),
	.cin(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~3 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N0
cycloneive_lcell_comb \ShiftLeft0~6 (
// Equation(s):
// \ShiftLeft0~6_combout  = (\ShiftLeft0~5_combout ) # ((\ShiftLeft0~4_combout ) # ((\ShiftLeft0~2_combout ) # (\ShiftLeft0~3_combout )))

	.dataa(\ShiftLeft0~5_combout ),
	.datab(\ShiftLeft0~4_combout ),
	.datac(\ShiftLeft0~2_combout ),
	.datad(\ShiftLeft0~3_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~6 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N16
cycloneive_lcell_comb \ShiftLeft0~7 (
// Equation(s):
// \ShiftLeft0~7_combout  = (Mux161) # ((\ShiftLeft0~6_combout ) # (Mux19))

	.dataa(gnd),
	.datab(Mux161),
	.datac(\ShiftLeft0~6_combout ),
	.datad(Mux19),
	.cin(gnd),
	.combout(\ShiftLeft0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~7 .lut_mask = 16'hFFFC;
defparam \ShiftLeft0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N10
cycloneive_lcell_comb \ShiftLeft0~11 (
// Equation(s):
// \ShiftLeft0~11_combout  = (\ShiftLeft0~8_combout ) # ((\ShiftLeft0~10_combout ) # (\ShiftLeft0~7_combout ))

	.dataa(\ShiftLeft0~8_combout ),
	.datab(\ShiftLeft0~10_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~7_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~11 .lut_mask = 16'hFFEE;
defparam \ShiftLeft0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N20
cycloneive_lcell_comb \Mux29~8 (
// Equation(s):
// \Mux29~8_combout  = (\Mux19~1_combout  & (((\Mux19~2_combout ) # (!\ShiftLeft0~11_combout )) # (!\Mux29~3_combout )))

	.dataa(\Mux19~1_combout ),
	.datab(\Mux29~3_combout ),
	.datac(\Mux19~2_combout ),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\Mux29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~8 .lut_mask = 16'hA2AA;
defparam \Mux29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N6
cycloneive_lcell_comb \Mux29~9 (
// Equation(s):
// \Mux29~9_combout  = (\Mux19~2_combout  & ((\Add0~13_combout ) # ((!\Mux29~8_combout )))) # (!\Mux19~2_combout  & (((\Mux29~7_combout  & \Mux29~8_combout ))))

	.dataa(\Add0~13_combout ),
	.datab(\Mux29~7_combout ),
	.datac(\Mux19~2_combout ),
	.datad(\Mux29~8_combout ),
	.cin(gnd),
	.combout(\Mux29~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~9 .lut_mask = 16'hACF0;
defparam \Mux29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N28
cycloneive_lcell_comb \Mux29~10 (
// Equation(s):
// \Mux29~10_combout  = (\Mux19~1_combout  & (((\Mux29~9_combout )))) # (!\Mux19~1_combout  & ((Mux291 & (!alu_a_mux_output_2 & !\Mux29~9_combout )) # (!Mux291 & (alu_a_mux_output_2 $ (\Mux29~9_combout )))))

	.dataa(\Mux19~1_combout ),
	.datab(Mux291),
	.datac(alu_a_mux_output_2),
	.datad(\Mux29~9_combout ),
	.cin(gnd),
	.combout(\Mux29~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~10 .lut_mask = 16'hAB14;
defparam \Mux29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N14
cycloneive_lcell_comb \ShiftRight0~37 (
// Equation(s):
// \ShiftRight0~37_combout  = (Mux301 & (alu_a_mux_output_14)) # (!Mux301 & ((alu_a_mux_output_12)))

	.dataa(Mux301),
	.datab(alu_a_mux_output_14),
	.datac(gnd),
	.datad(alu_a_mux_output_12),
	.cin(gnd),
	.combout(\ShiftRight0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~37 .lut_mask = 16'hDD88;
defparam \ShiftRight0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N0
cycloneive_lcell_comb \ShiftRight0~60 (
// Equation(s):
// \ShiftRight0~60_combout  = (Mux301 & (alu_a_mux_output_13)) # (!Mux301 & ((alu_a_mux_output_11)))

	.dataa(alu_a_mux_output_13),
	.datab(gnd),
	.datac(alu_a_mux_output_11),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftRight0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~60 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N28
cycloneive_lcell_comb \ShiftRight0~76 (
// Equation(s):
// \ShiftRight0~76_combout  = (Mux311 & (\ShiftRight0~37_combout )) # (!Mux311 & ((\ShiftRight0~60_combout )))

	.dataa(gnd),
	.datab(Mux311),
	.datac(\ShiftRight0~37_combout ),
	.datad(\ShiftRight0~60_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~76 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y40_N16
cycloneive_lcell_comb \ShiftRight0~77 (
// Equation(s):
// \ShiftRight0~77_combout  = (!Mux301 & ((Mux311 & (alu_a_mux_output_16)) # (!Mux311 & ((alu_a_mux_output_15)))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_16),
	.datac(alu_a_mux_output_15),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftRight0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~77 .lut_mask = 16'h4450;
defparam \ShiftRight0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y40_N14
cycloneive_lcell_comb \ShiftRight0~78 (
// Equation(s):
// \ShiftRight0~78_combout  = (Mux301 & ((Mux311 & (alu_a_mux_output_18)) # (!Mux311 & ((alu_a_mux_output_17)))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_18),
	.datac(alu_a_mux_output_17),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftRight0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~78 .lut_mask = 16'h88A0;
defparam \ShiftRight0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N8
cycloneive_lcell_comb \ShiftRight0~79 (
// Equation(s):
// \ShiftRight0~79_combout  = (Mux291 & (((\ShiftRight0~77_combout ) # (\ShiftRight0~78_combout )))) # (!Mux291 & (\ShiftRight0~76_combout ))

	.dataa(Mux291),
	.datab(\ShiftRight0~76_combout ),
	.datac(\ShiftRight0~77_combout ),
	.datad(\ShiftRight0~78_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~79 .lut_mask = 16'hEEE4;
defparam \ShiftRight0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N2
cycloneive_lcell_comb \ShiftRight0~6 (
// Equation(s):
// \ShiftRight0~6_combout  = (Mux311 & ((alu_a_mux_output_6))) # (!Mux311 & (alu_a_mux_output_5))

	.dataa(Mux311),
	.datab(alu_a_mux_output_5),
	.datac(gnd),
	.datad(alu_a_mux_output_6),
	.cin(gnd),
	.combout(\ShiftRight0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~6 .lut_mask = 16'hEE44;
defparam \ShiftRight0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N22
cycloneive_lcell_comb \ShiftRight0~59 (
// Equation(s):
// \ShiftRight0~59_combout  = (!Mux291 & !Mux281)

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux291),
	.datad(Mux281),
	.cin(gnd),
	.combout(\ShiftRight0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~59 .lut_mask = 16'h000F;
defparam \ShiftRight0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N30
cycloneive_lcell_comb \ShiftRight0~39 (
// Equation(s):
// \ShiftRight0~39_combout  = (Mux301 & ((alu_a_mux_output_10))) # (!Mux301 & (alu_a_mux_output_8))

	.dataa(alu_a_mux_output_8),
	.datab(gnd),
	.datac(alu_a_mux_output_10),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftRight0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~39 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N6
cycloneive_lcell_comb \ShiftRight0~75 (
// Equation(s):
// \ShiftRight0~75_combout  = (Mux311 & ((\ShiftRight0~39_combout ))) # (!Mux311 & (\ShiftRight0~57_combout ))

	.dataa(Mux311),
	.datab(gnd),
	.datac(\ShiftRight0~57_combout ),
	.datad(\ShiftRight0~39_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~75 .lut_mask = 16'hFA50;
defparam \ShiftRight0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N28
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (\ShiftRight0~59_combout  & (\ShiftRight0~3_combout  & (!\Mux29~0_combout ))) # (!\ShiftRight0~59_combout  & (((\Mux29~0_combout ) # (\ShiftRight0~75_combout ))))

	.dataa(\ShiftRight0~3_combout ),
	.datab(\ShiftRight0~59_combout ),
	.datac(\Mux29~0_combout ),
	.datad(\ShiftRight0~75_combout ),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'h3B38;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N14
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (\Mux29~0_combout  & ((\Mux28~0_combout  & (\ShiftRight0~79_combout )) # (!\Mux28~0_combout  & ((\ShiftRight0~6_combout ))))) # (!\Mux29~0_combout  & (((\Mux28~0_combout ))))

	.dataa(\Mux29~0_combout ),
	.datab(\ShiftRight0~79_combout ),
	.datac(\ShiftRight0~6_combout ),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hDDA0;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N18
cycloneive_lcell_comb \Mux29~5 (
// Equation(s):
// \Mux29~5_combout  = (temp_ALUop_output_1) # ((temp_ALUop_output_0 & Mux271))

	.dataa(temp_ALUop_output_0),
	.datab(temp_ALUop_output_1),
	.datac(gnd),
	.datad(Mux271),
	.cin(gnd),
	.combout(\Mux29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~5 .lut_mask = 16'hEECC;
defparam \Mux29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N20
cycloneive_lcell_comb \ShiftLeft0~20 (
// Equation(s):
// \ShiftLeft0~20_combout  = (!Mux301 & ((Mux311 & (alu_a_mux_output_2)) # (!Mux311 & ((alu_a_mux_output_31)))))

	.dataa(alu_a_mux_output_2),
	.datab(Mux311),
	.datac(alu_a_mux_output_31),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftLeft0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~20 .lut_mask = 16'h00B8;
defparam \ShiftLeft0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N26
cycloneive_lcell_comb \ShiftLeft0~21 (
// Equation(s):
// \ShiftLeft0~21_combout  = (\ShiftRight0~59_combout  & ((\ShiftLeft0~20_combout ) # ((\ShiftLeft0~12_combout  & Mux301))))

	.dataa(\ShiftLeft0~12_combout ),
	.datab(\ShiftRight0~59_combout ),
	.datac(Mux301),
	.datad(\ShiftLeft0~20_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~21 .lut_mask = 16'hCC80;
defparam \ShiftLeft0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N4
cycloneive_lcell_comb \ShiftLeft0~8 (
// Equation(s):
// \ShiftLeft0~8_combout  = (Mux21) # ((Mux17) # ((!Mux16 & alu_b_mux_output_14)))

	.dataa(Mux16),
	.datab(Mux21),
	.datac(alu_b_mux_output_14),
	.datad(Mux17),
	.cin(gnd),
	.combout(\ShiftLeft0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~8 .lut_mask = 16'hFFDC;
defparam \ShiftLeft0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N0
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (!Mux271 & (!\ShiftLeft0~7_combout  & (!\ShiftLeft0~10_combout  & !\ShiftLeft0~8_combout )))

	.dataa(Mux271),
	.datab(\ShiftLeft0~7_combout ),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\ShiftLeft0~8_combout ),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'h0001;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N10
cycloneive_lcell_comb \Mux29~4 (
// Equation(s):
// \Mux29~4_combout  = (temp_ALUop_output_1) # ((!temp_ALUop_output_0 & \Mux19~0_combout ))

	.dataa(temp_ALUop_output_0),
	.datab(gnd),
	.datac(\Mux19~0_combout ),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Mux29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~4 .lut_mask = 16'hFF50;
defparam \Mux29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N20
cycloneive_lcell_comb \Mux28~2 (
// Equation(s):
// \Mux28~2_combout  = (\Mux29~5_combout  & ((\OUTPUT~1_combout ) # ((!\Mux29~4_combout )))) # (!\Mux29~5_combout  & (((\ShiftLeft0~21_combout  & \Mux29~4_combout ))))

	.dataa(\OUTPUT~1_combout ),
	.datab(\Mux29~5_combout ),
	.datac(\ShiftLeft0~21_combout ),
	.datad(\Mux29~4_combout ),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~2 .lut_mask = 16'hB8CC;
defparam \Mux28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N16
cycloneive_lcell_comb \Mux28~3 (
// Equation(s):
// \Mux28~3_combout  = (\Mux29~3_combout  & ((\Mux28~2_combout  & (\ShiftRight0~89_combout )) # (!\Mux28~2_combout  & ((\Mux28~1_combout ))))) # (!\Mux29~3_combout  & (((\Mux28~2_combout ))))

	.dataa(\ShiftRight0~89_combout ),
	.datab(\Mux28~1_combout ),
	.datac(\Mux29~3_combout ),
	.datad(\Mux28~2_combout ),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~3 .lut_mask = 16'hAFC0;
defparam \Mux28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N22
cycloneive_lcell_comb \Mux28~4 (
// Equation(s):
// \Mux28~4_combout  = (\Mux29~8_combout  & ((\Mux19~2_combout  & (\Add0~16_combout )) # (!\Mux19~2_combout  & ((\Mux28~3_combout ))))) # (!\Mux29~8_combout  & (((\Mux19~2_combout ))))

	.dataa(\Add0~16_combout ),
	.datab(\Mux29~8_combout ),
	.datac(\Mux19~2_combout ),
	.datad(\Mux28~3_combout ),
	.cin(gnd),
	.combout(\Mux28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~4 .lut_mask = 16'hBCB0;
defparam \Mux28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N6
cycloneive_lcell_comb \Mux28~5 (
// Equation(s):
// \Mux28~5_combout  = (\Mux28~4_combout  & ((\Mux19~1_combout ) # ((!Mux281 & !alu_a_mux_output_31)))) # (!\Mux28~4_combout  & (!\Mux19~1_combout  & (Mux281 $ (alu_a_mux_output_31))))

	.dataa(Mux281),
	.datab(alu_a_mux_output_31),
	.datac(\Mux28~4_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~5 .lut_mask = 16'hF016;
defparam \Mux28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N18
cycloneive_lcell_comb \Mux26~5 (
// Equation(s):
// \Mux26~5_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!alu_a_mux_output_5 & !Mux26)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (alu_a_mux_output_5 $ (Mux26))))

	.dataa(alu_a_mux_output_5),
	.datab(Mux26),
	.datac(\Mux19~2_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~5 .lut_mask = 16'hF016;
defparam \Mux26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N18
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = temp_ALUop_output_0 $ (((temp_ALUsrc_output_0 & ((temp_imemload_output_5) # (temp_ALUsrc_output_1))) # (!temp_ALUsrc_output_0 & ((!temp_ALUsrc_output_1)))))

	.dataa(temp_ALUop_output_0),
	.datab(temp_imemload_output_5),
	.datac(temp_ALUsrc_output_0),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(\Add0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h5A65;
defparam \Add0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N8
cycloneive_lcell_comb \Add0~19 (
// Equation(s):
// \Add0~19_combout  = \Add0~18_combout  $ (((!alu_b_mux_output_5 & (temp_ALUsrc_output_1 $ (!temp_ALUsrc_output_0)))))

	.dataa(temp_ALUsrc_output_1),
	.datab(\Add0~18_combout ),
	.datac(temp_ALUsrc_output_0),
	.datad(alu_b_mux_output_5),
	.cin(gnd),
	.combout(\Add0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~19 .lut_mask = 16'hCC69;
defparam \Add0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N10
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = temp_ALUop_output_0 $ (((Mux27) # ((!Mux16 & alu_b_mux_output_4))))

	.dataa(temp_ALUop_output_0),
	.datab(Mux16),
	.datac(Mux27),
	.datad(alu_b_mux_output_4),
	.cin(gnd),
	.combout(\Add0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'h595A;
defparam \Add0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N16
cycloneive_lcell_comb \Add0~15 (
// Equation(s):
// \Add0~15_combout  = temp_ALUop_output_0 $ (((Mux28) # ((!Mux16 & alu_b_mux_output_3))))

	.dataa(temp_ALUop_output_0),
	.datab(Mux16),
	.datac(Mux28),
	.datad(alu_b_mux_output_3),
	.cin(gnd),
	.combout(\Add0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~15 .lut_mask = 16'h595A;
defparam \Add0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N24
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = temp_ALUop_output_0 $ (((Mux29) # ((!Mux16 & alu_b_mux_output_2))))

	.dataa(temp_ALUop_output_0),
	.datab(Mux16),
	.datac(Mux29),
	.datad(alu_b_mux_output_2),
	.cin(gnd),
	.combout(\Add0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'h595A;
defparam \Add0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N26
cycloneive_lcell_comb \Add0~21 (
// Equation(s):
// \Add0~21_combout  = (alu_a_mux_output_4 & ((\Add0~20_combout  & (\Add0~17  & VCC)) # (!\Add0~20_combout  & (!\Add0~17 )))) # (!alu_a_mux_output_4 & ((\Add0~20_combout  & (!\Add0~17 )) # (!\Add0~20_combout  & ((\Add0~17 ) # (GND)))))
// \Add0~22  = CARRY((alu_a_mux_output_4 & (!\Add0~20_combout  & !\Add0~17 )) # (!alu_a_mux_output_4 & ((!\Add0~17 ) # (!\Add0~20_combout ))))

	.dataa(alu_a_mux_output_4),
	.datab(\Add0~20_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~21_combout ),
	.cout(\Add0~22 ));
// synopsys translate_off
defparam \Add0~21 .lut_mask = 16'h9617;
defparam \Add0~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N28
cycloneive_lcell_comb \Add0~23 (
// Equation(s):
// \Add0~23_combout  = ((alu_a_mux_output_5 $ (\Add0~19_combout  $ (!\Add0~22 )))) # (GND)
// \Add0~24  = CARRY((alu_a_mux_output_5 & ((\Add0~19_combout ) # (!\Add0~22 ))) # (!alu_a_mux_output_5 & (\Add0~19_combout  & !\Add0~22 )))

	.dataa(alu_a_mux_output_5),
	.datab(\Add0~19_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~22 ),
	.combout(\Add0~23_combout ),
	.cout(\Add0~24 ));
// synopsys translate_off
defparam \Add0~23 .lut_mask = 16'h698E;
defparam \Add0~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N2
cycloneive_lcell_comb \Mux27~3 (
// Equation(s):
// \Mux27~3_combout  = (Mux281) # (Mux271)

	.dataa(Mux281),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux271),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~3 .lut_mask = 16'hFFAA;
defparam \Mux27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N24
cycloneive_lcell_comb \Mux27~2 (
// Equation(s):
// \Mux27~2_combout  = (Mux271) # ((Mux291 & !Mux281))

	.dataa(gnd),
	.datab(Mux291),
	.datac(Mux281),
	.datad(Mux271),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~2 .lut_mask = 16'hFF0C;
defparam \Mux27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N4
cycloneive_lcell_comb \ShiftRight0~23 (
// Equation(s):
// \ShiftRight0~23_combout  = (Mux301 & ((Mux311 & (alu_a_mux_output_20)) # (!Mux311 & ((alu_a_mux_output_19)))))

	.dataa(alu_a_mux_output_20),
	.datab(Mux311),
	.datac(Mux301),
	.datad(alu_a_mux_output_19),
	.cin(gnd),
	.combout(\ShiftRight0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~23 .lut_mask = 16'hB080;
defparam \ShiftRight0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N10
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (!Mux301 & Mux311)

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux301),
	.datad(Mux311),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'h0F00;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N12
cycloneive_lcell_comb \ShiftRight0~24 (
// Equation(s):
// \ShiftRight0~24_combout  = (\ShiftRight0~22_combout ) # ((\ShiftRight0~23_combout ) # ((alu_a_mux_output_18 & \Mux1~0_combout )))

	.dataa(\ShiftRight0~22_combout ),
	.datab(\ShiftRight0~23_combout ),
	.datac(alu_a_mux_output_18),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~24 .lut_mask = 16'hFEEE;
defparam \ShiftRight0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N26
cycloneive_lcell_comb \ShiftRight0~10 (
// Equation(s):
// \ShiftRight0~10_combout  = (Mux301 & (alu_a_mux_output_15)) # (!Mux301 & ((alu_a_mux_output_13)))

	.dataa(gnd),
	.datab(alu_a_mux_output_15),
	.datac(alu_a_mux_output_13),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftRight0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~10 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N24
cycloneive_lcell_comb \ShiftRight0~9 (
// Equation(s):
// \ShiftRight0~9_combout  = (Mux311 & ((Mux301 & ((alu_a_mux_output_16))) # (!Mux301 & (alu_a_mux_output_14))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_14),
	.datac(Mux311),
	.datad(alu_a_mux_output_16),
	.cin(gnd),
	.combout(\ShiftRight0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~9 .lut_mask = 16'hE040;
defparam \ShiftRight0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N28
cycloneive_lcell_comb \ShiftRight0~11 (
// Equation(s):
// \ShiftRight0~11_combout  = (\ShiftRight0~9_combout ) # ((!Mux311 & \ShiftRight0~10_combout ))

	.dataa(gnd),
	.datab(Mux311),
	.datac(\ShiftRight0~10_combout ),
	.datad(\ShiftRight0~9_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~11 .lut_mask = 16'hFF30;
defparam \ShiftRight0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N4
cycloneive_lcell_comb \ShiftRight0~90 (
// Equation(s):
// \ShiftRight0~90_combout  = (Mux291 & (\ShiftRight0~24_combout )) # (!Mux291 & ((\ShiftRight0~11_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~24_combout ),
	.datac(Mux291),
	.datad(\ShiftRight0~11_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~90 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N20
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (\Mux27~3_combout  & (((\Mux27~2_combout ) # (\ShiftRight0~90_combout )))) # (!\Mux27~3_combout  & (\ShiftRight0~7_combout  & (!\Mux27~2_combout )))

	.dataa(\ShiftRight0~7_combout ),
	.datab(\Mux27~3_combout ),
	.datac(\Mux27~2_combout ),
	.datad(\ShiftRight0~90_combout ),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hCEC2;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N28
cycloneive_lcell_comb \ShiftRight0~19 (
// Equation(s):
// \ShiftRight0~19_combout  = (Mux301 & ((Mux311 & (alu_a_mux_output_28)) # (!Mux311 & ((alu_a_mux_output_27))))) # (!Mux301 & (((Mux311))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_28),
	.datac(Mux311),
	.datad(alu_a_mux_output_27),
	.cin(gnd),
	.combout(\ShiftRight0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~19 .lut_mask = 16'hDAD0;
defparam \ShiftRight0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N30
cycloneive_lcell_comb \ShiftRight0~20 (
// Equation(s):
// \ShiftRight0~20_combout  = (Mux301 & (((\ShiftRight0~19_combout )))) # (!Mux301 & ((\ShiftRight0~19_combout  & ((alu_a_mux_output_26))) # (!\ShiftRight0~19_combout  & (alu_a_mux_output_25))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_25),
	.datac(alu_a_mux_output_26),
	.datad(\ShiftRight0~19_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~20 .lut_mask = 16'hFA44;
defparam \ShiftRight0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N12
cycloneive_lcell_comb \ShiftRight0~26 (
// Equation(s):
// \ShiftRight0~26_combout  = (!Mux301 & ((Mux311 & ((alu_a_mux_output_22))) # (!Mux311 & (alu_a_mux_output_21))))

	.dataa(alu_a_mux_output_21),
	.datab(Mux301),
	.datac(Mux311),
	.datad(alu_a_mux_output_22),
	.cin(gnd),
	.combout(\ShiftRight0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~26 .lut_mask = 16'h3202;
defparam \ShiftRight0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N2
cycloneive_lcell_comb \ShiftRight0~91 (
// Equation(s):
// \ShiftRight0~91_combout  = (Mux291 & (((\ShiftRight0~20_combout )))) # (!Mux291 & ((\ShiftRight0~25_combout ) # ((\ShiftRight0~26_combout ))))

	.dataa(\ShiftRight0~25_combout ),
	.datab(\ShiftRight0~20_combout ),
	.datac(\ShiftRight0~26_combout ),
	.datad(Mux291),
	.cin(gnd),
	.combout(\ShiftRight0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~91 .lut_mask = 16'hCCFA;
defparam \ShiftRight0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N16
cycloneive_lcell_comb \ShiftRight0~92 (
// Equation(s):
// \ShiftRight0~92_combout  = (Mux281 & (\ShiftRight0~18_combout  & (!Mux291))) # (!Mux281 & (((\ShiftRight0~91_combout ))))

	.dataa(\ShiftRight0~18_combout ),
	.datab(Mux281),
	.datac(Mux291),
	.datad(\ShiftRight0~91_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~92 .lut_mask = 16'h3B08;
defparam \ShiftRight0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N16
cycloneive_lcell_comb \ShiftRight0~12 (
// Equation(s):
// \ShiftRight0~12_combout  = (Mux301 & ((alu_a_mux_output_12))) # (!Mux301 & (alu_a_mux_output_10))

	.dataa(Mux301),
	.datab(gnd),
	.datac(alu_a_mux_output_10),
	.datad(alu_a_mux_output_12),
	.cin(gnd),
	.combout(\ShiftRight0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~12 .lut_mask = 16'hFA50;
defparam \ShiftRight0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N2
cycloneive_lcell_comb \ShiftRight0~13 (
// Equation(s):
// \ShiftRight0~13_combout  = (Mux301 & (alu_a_mux_output_11)) # (!Mux301 & ((alu_a_mux_output_9)))

	.dataa(gnd),
	.datab(alu_a_mux_output_11),
	.datac(alu_a_mux_output_9),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftRight0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~13 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N4
cycloneive_lcell_comb \ShiftRight0~14 (
// Equation(s):
// \ShiftRight0~14_combout  = (Mux311 & (\ShiftRight0~12_combout )) # (!Mux311 & ((\ShiftRight0~13_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~12_combout ),
	.datac(Mux311),
	.datad(\ShiftRight0~13_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~14 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N10
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (\Mux27~2_combout  & ((\Mux26~0_combout  & (\ShiftRight0~92_combout )) # (!\Mux26~0_combout  & ((\ShiftRight0~14_combout ))))) # (!\Mux27~2_combout  & (\Mux26~0_combout ))

	.dataa(\Mux27~2_combout ),
	.datab(\Mux26~0_combout ),
	.datac(\ShiftRight0~92_combout ),
	.datad(\ShiftRight0~14_combout ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hE6C4;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N22
cycloneive_lcell_comb \ShiftLeft0~26 (
// Equation(s):
// \ShiftLeft0~26_combout  = (\ShiftLeft0~8_combout ) # ((\ShiftLeft0~6_combout ) # ((Mux161) # (Mux19)))

	.dataa(\ShiftLeft0~8_combout ),
	.datab(\ShiftLeft0~6_combout ),
	.datac(Mux161),
	.datad(Mux19),
	.cin(gnd),
	.combout(\ShiftLeft0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~26 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N12
cycloneive_lcell_comb \Mux27~4 (
// Equation(s):
// \Mux27~4_combout  = (!temp_ALUop_output_1 & (((!\ShiftLeft0~10_combout  & !\ShiftLeft0~26_combout )) # (!temp_ALUop_output_0)))

	.dataa(temp_ALUop_output_1),
	.datab(\ShiftLeft0~10_combout ),
	.datac(temp_ALUop_output_0),
	.datad(\ShiftLeft0~26_combout ),
	.cin(gnd),
	.combout(\Mux27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~4 .lut_mask = 16'h0515;
defparam \Mux27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N8
cycloneive_lcell_comb \Mux26~3 (
// Equation(s):
// \Mux26~3_combout  = (temp_ALUop_output_0 & (((\Mux26~1_combout  & \Mux27~4_combout )))) # (!temp_ALUop_output_0 & ((\Mux26~2_combout ) # ((!\Mux27~4_combout ))))

	.dataa(\Mux26~2_combout ),
	.datab(\Mux26~1_combout ),
	.datac(temp_ALUop_output_0),
	.datad(\Mux27~4_combout ),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~3 .lut_mask = 16'hCA0F;
defparam \Mux26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N2
cycloneive_lcell_comb \Mux26~4 (
// Equation(s):
// \Mux26~4_combout  = (\Mux26~3_combout  & (((alu_a_mux_output_5 & Mux26)) # (!temp_ALUop_output_1))) # (!\Mux26~3_combout  & (temp_ALUop_output_1 & ((alu_a_mux_output_5) # (Mux26))))

	.dataa(alu_a_mux_output_5),
	.datab(Mux26),
	.datac(\Mux26~3_combout ),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Mux26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~4 .lut_mask = 16'h8EF0;
defparam \Mux26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N14
cycloneive_lcell_comb \Mux27~12 (
// Equation(s):
// \Mux27~12_combout  = (Mux27) # ((alu_b_mux_output_4 & (temp_ALUsrc_output_0 $ (!temp_ALUsrc_output_1))))

	.dataa(temp_ALUsrc_output_0),
	.datab(temp_ALUsrc_output_1),
	.datac(Mux27),
	.datad(alu_b_mux_output_4),
	.cin(gnd),
	.combout(\Mux27~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~12 .lut_mask = 16'hF9F0;
defparam \Mux27~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N6
cycloneive_lcell_comb \Mux27~10 (
// Equation(s):
// \Mux27~10_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!\Mux27~12_combout  & !alu_a_mux_output_4)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (\Mux27~12_combout  $ (alu_a_mux_output_4))))

	.dataa(\Mux27~12_combout ),
	.datab(alu_a_mux_output_4),
	.datac(\Mux19~2_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux27~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~10 .lut_mask = 16'hF016;
defparam \Mux27~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N20
cycloneive_lcell_comb \ShiftRight0~53 (
// Equation(s):
// \ShiftRight0~53_combout  = (Mux301 & ((Mux311 & ((alu_a_mux_output_27))) # (!Mux311 & (alu_a_mux_output_26)))) # (!Mux301 & (Mux311))

	.dataa(Mux301),
	.datab(Mux311),
	.datac(alu_a_mux_output_26),
	.datad(alu_a_mux_output_27),
	.cin(gnd),
	.combout(\ShiftRight0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~53 .lut_mask = 16'hEC64;
defparam \ShiftRight0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N14
cycloneive_lcell_comb \ShiftRight0~54 (
// Equation(s):
// \ShiftRight0~54_combout  = (Mux301 & (((\ShiftRight0~53_combout )))) # (!Mux301 & ((\ShiftRight0~53_combout  & ((alu_a_mux_output_25))) # (!\ShiftRight0~53_combout  & (alu_a_mux_output_24))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_24),
	.datac(alu_a_mux_output_25),
	.datad(\ShiftRight0~53_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~54 .lut_mask = 16'hFA44;
defparam \ShiftRight0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N30
cycloneive_lcell_comb \ShiftRight0~46 (
// Equation(s):
// \ShiftRight0~46_combout  = (!Mux301 & ((Mux311 & (alu_a_mux_output_21)) # (!Mux311 & ((alu_a_mux_output_20)))))

	.dataa(alu_a_mux_output_21),
	.datab(Mux311),
	.datac(Mux301),
	.datad(alu_a_mux_output_20),
	.cin(gnd),
	.combout(\ShiftRight0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~46 .lut_mask = 16'h0B08;
defparam \ShiftRight0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N16
cycloneive_lcell_comb \ShiftRight0~94 (
// Equation(s):
// \ShiftRight0~94_combout  = (Mux291 & (((\ShiftRight0~54_combout )))) # (!Mux291 & ((\ShiftRight0~47_combout ) # ((\ShiftRight0~46_combout ))))

	.dataa(\ShiftRight0~47_combout ),
	.datab(\ShiftRight0~54_combout ),
	.datac(Mux291),
	.datad(\ShiftRight0~46_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~94 .lut_mask = 16'hCFCA;
defparam \ShiftRight0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N8
cycloneive_lcell_comb \ShiftRight0~43 (
// Equation(s):
// \ShiftRight0~43_combout  = (!Mux301 & ((Mux311 & ((alu_a_mux_output_29))) # (!Mux311 & (alu_a_mux_output_28))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_28),
	.datac(Mux311),
	.datad(alu_a_mux_output_29),
	.cin(gnd),
	.combout(\ShiftRight0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~43 .lut_mask = 16'h5404;
defparam \ShiftRight0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N6
cycloneive_lcell_comb \ShiftRight0~45 (
// Equation(s):
// \ShiftRight0~45_combout  = (\ShiftRight0~43_combout ) # ((Mux301 & \ShiftRight0~44_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~43_combout ),
	.datac(Mux301),
	.datad(\ShiftRight0~44_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~45 .lut_mask = 16'hFCCC;
defparam \ShiftRight0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N10
cycloneive_lcell_comb \ShiftRight0~95 (
// Equation(s):
// \ShiftRight0~95_combout  = (Mux281 & (((!Mux291 & \ShiftRight0~45_combout )))) # (!Mux281 & (\ShiftRight0~94_combout ))

	.dataa(Mux281),
	.datab(\ShiftRight0~94_combout ),
	.datac(Mux291),
	.datad(\ShiftRight0~45_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~95 .lut_mask = 16'h4E44;
defparam \ShiftRight0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N0
cycloneive_lcell_comb \ShiftRight0~40 (
// Equation(s):
// \ShiftRight0~40_combout  = (Mux311 & ((\ShiftRight0~13_combout ))) # (!Mux311 & (\ShiftRight0~39_combout ))

	.dataa(gnd),
	.datab(Mux311),
	.datac(\ShiftRight0~39_combout ),
	.datad(\ShiftRight0~13_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~40 .lut_mask = 16'hFC30;
defparam \ShiftRight0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N14
cycloneive_lcell_comb \ShiftRight0~33 (
// Equation(s):
// \ShiftRight0~33_combout  = (Mux301 & ((Mux311 & (alu_a_mux_output_7)) # (!Mux311 & ((alu_a_mux_output_6)))))

	.dataa(Mux311),
	.datab(Mux301),
	.datac(alu_a_mux_output_7),
	.datad(alu_a_mux_output_6),
	.cin(gnd),
	.combout(\ShiftRight0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~33 .lut_mask = 16'hC480;
defparam \ShiftRight0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N10
cycloneive_lcell_comb \ShiftRight0~35 (
// Equation(s):
// \ShiftRight0~35_combout  = (\ShiftRight0~33_combout ) # ((!Mux301 & \ShiftRight0~34_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~33_combout ),
	.datac(Mux301),
	.datad(\ShiftRight0~34_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~35 .lut_mask = 16'hCFCC;
defparam \ShiftRight0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N4
cycloneive_lcell_comb \Mux27~5 (
// Equation(s):
// \Mux27~5_combout  = (\Mux27~3_combout  & (\Mux27~2_combout )) # (!\Mux27~3_combout  & ((\Mux27~2_combout  & (\ShiftRight0~40_combout )) # (!\Mux27~2_combout  & ((\ShiftRight0~35_combout )))))

	.dataa(\Mux27~3_combout ),
	.datab(\Mux27~2_combout ),
	.datac(\ShiftRight0~40_combout ),
	.datad(\ShiftRight0~35_combout ),
	.cin(gnd),
	.combout(\Mux27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~5 .lut_mask = 16'hD9C8;
defparam \Mux27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N2
cycloneive_lcell_comb \Mux27~6 (
// Equation(s):
// \Mux27~6_combout  = (\Mux27~5_combout  & (((\ShiftRight0~95_combout ) # (!\Mux27~3_combout )))) # (!\Mux27~5_combout  & (\ShiftRight0~93_combout  & ((\Mux27~3_combout ))))

	.dataa(\ShiftRight0~93_combout ),
	.datab(\ShiftRight0~95_combout ),
	.datac(\Mux27~5_combout ),
	.datad(\Mux27~3_combout ),
	.cin(gnd),
	.combout(\Mux27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~6 .lut_mask = 16'hCAF0;
defparam \Mux27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N18
cycloneive_lcell_comb \ShiftLeft0~22 (
// Equation(s):
// \ShiftLeft0~22_combout  = (Mux301 & ((alu_a_mux_output_2))) # (!Mux301 & (alu_a_mux_output_4))

	.dataa(Mux301),
	.datab(gnd),
	.datac(alu_a_mux_output_4),
	.datad(alu_a_mux_output_2),
	.cin(gnd),
	.combout(\ShiftLeft0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~22 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N0
cycloneive_lcell_comb \ShiftLeft0~28 (
// Equation(s):
// \ShiftLeft0~28_combout  = (Mux311 & (\ShiftLeft0~27_combout )) # (!Mux311 & ((\ShiftLeft0~22_combout )))

	.dataa(\ShiftLeft0~27_combout ),
	.datab(\ShiftLeft0~22_combout ),
	.datac(gnd),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftLeft0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~28 .lut_mask = 16'hAACC;
defparam \ShiftLeft0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N0
cycloneive_lcell_comb \ShiftLeft0~16 (
// Equation(s):
// \ShiftLeft0~16_combout  = (!Mux301 & (alu_a_mux_output_0 & !Mux311))

	.dataa(Mux301),
	.datab(gnd),
	.datac(alu_a_mux_output_0),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftLeft0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~16 .lut_mask = 16'h0050;
defparam \ShiftLeft0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N12
cycloneive_lcell_comb \ShiftLeft0~29 (
// Equation(s):
// \ShiftLeft0~29_combout  = (Mux291 & ((\ShiftLeft0~16_combout ))) # (!Mux291 & (\ShiftLeft0~28_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~28_combout ),
	.datac(Mux291),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~29 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N6
cycloneive_lcell_comb \Mux27~7 (
// Equation(s):
// \Mux27~7_combout  = (!Mux281 & (\ShiftLeft0~29_combout  & \Mux19~0_combout ))

	.dataa(Mux281),
	.datab(\ShiftLeft0~29_combout ),
	.datac(\Mux19~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~7 .lut_mask = 16'h4040;
defparam \Mux27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N16
cycloneive_lcell_comb \Mux27~8 (
// Equation(s):
// \Mux27~8_combout  = (\Mux27~4_combout  & ((temp_ALUop_output_0 & (\Mux27~6_combout )) # (!temp_ALUop_output_0 & ((\Mux27~7_combout ))))) # (!\Mux27~4_combout  & (((!temp_ALUop_output_0))))

	.dataa(\Mux27~4_combout ),
	.datab(\Mux27~6_combout ),
	.datac(temp_ALUop_output_0),
	.datad(\Mux27~7_combout ),
	.cin(gnd),
	.combout(\Mux27~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~8 .lut_mask = 16'h8F85;
defparam \Mux27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N16
cycloneive_lcell_comb \Mux27~9 (
// Equation(s):
// \Mux27~9_combout  = (temp_ALUop_output_1 & ((alu_a_mux_output_4 & ((Mux271) # (!\Mux27~8_combout ))) # (!alu_a_mux_output_4 & (Mux271 & !\Mux27~8_combout )))) # (!temp_ALUop_output_1 & (((\Mux27~8_combout ))))

	.dataa(alu_a_mux_output_4),
	.datab(temp_ALUop_output_1),
	.datac(Mux271),
	.datad(\Mux27~8_combout ),
	.cin(gnd),
	.combout(\Mux27~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~9 .lut_mask = 16'hB3C8;
defparam \Mux27~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N10
cycloneive_lcell_comb \Mux24~5 (
// Equation(s):
// \Mux24~5_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!alu_a_mux_output_7 & !Mux24)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (alu_a_mux_output_7 $ (Mux24))))

	.dataa(\Mux19~2_combout ),
	.datab(alu_a_mux_output_7),
	.datac(Mux24),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~5 .lut_mask = 16'hAA16;
defparam \Mux24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N2
cycloneive_lcell_comb \ShiftRight0~80 (
// Equation(s):
// \ShiftRight0~80_combout  = (!Mux301 & (alu_a_mux_output_311 & !Mux311))

	.dataa(Mux301),
	.datab(gnd),
	.datac(alu_a_mux_output_311),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftRight0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~80 .lut_mask = 16'h0050;
defparam \ShiftRight0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N18
cycloneive_lcell_comb \ShiftRight0~82 (
// Equation(s):
// \ShiftRight0~82_combout  = (!Mux311 & ((Mux301 & (alu_a_mux_output_29)) # (!Mux301 & ((alu_a_mux_output_27)))))

	.dataa(alu_a_mux_output_29),
	.datab(Mux301),
	.datac(Mux311),
	.datad(alu_a_mux_output_27),
	.cin(gnd),
	.combout(\ShiftRight0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~82 .lut_mask = 16'h0B08;
defparam \ShiftRight0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N16
cycloneive_lcell_comb \ShiftRight0~81 (
// Equation(s):
// \ShiftRight0~81_combout  = (Mux311 & ((Mux301 & (alu_a_mux_output_30)) # (!Mux301 & ((alu_a_mux_output_28)))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_30),
	.datac(alu_a_mux_output_28),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftRight0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~81 .lut_mask = 16'hD800;
defparam \ShiftRight0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N12
cycloneive_lcell_comb \ShiftRight0~97 (
// Equation(s):
// \ShiftRight0~97_combout  = (Mux291 & (((\ShiftRight0~82_combout ) # (\ShiftRight0~81_combout )))) # (!Mux291 & (\ShiftRight0~85_combout ))

	.dataa(\ShiftRight0~85_combout ),
	.datab(\ShiftRight0~82_combout ),
	.datac(\ShiftRight0~81_combout ),
	.datad(Mux291),
	.cin(gnd),
	.combout(\ShiftRight0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~97 .lut_mask = 16'hFCAA;
defparam \ShiftRight0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N2
cycloneive_lcell_comb \ShiftRight0~98 (
// Equation(s):
// \ShiftRight0~98_combout  = (Mux281 & (!Mux291 & (\ShiftRight0~80_combout ))) # (!Mux281 & (((\ShiftRight0~97_combout ))))

	.dataa(Mux291),
	.datab(Mux281),
	.datac(\ShiftRight0~80_combout ),
	.datad(\ShiftRight0~97_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~98 .lut_mask = 16'h7340;
defparam \ShiftRight0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N0
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (\Mux24~0_combout  & (((\ShiftRight0~98_combout )) # (!\Mux27~2_combout ))) # (!\Mux24~0_combout  & (\Mux27~2_combout  & ((\ShiftRight0~76_combout ))))

	.dataa(\Mux24~0_combout ),
	.datab(\Mux27~2_combout ),
	.datac(\ShiftRight0~98_combout ),
	.datad(\ShiftRight0~76_combout ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hE6A2;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N22
cycloneive_lcell_comb \ShiftLeft0~32 (
// Equation(s):
// \ShiftLeft0~32_combout  = (Mux301 & ((alu_a_mux_output_5))) # (!Mux301 & (alu_a_mux_output_7))

	.dataa(gnd),
	.datab(Mux301),
	.datac(alu_a_mux_output_7),
	.datad(alu_a_mux_output_5),
	.cin(gnd),
	.combout(\ShiftLeft0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~32 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N16
cycloneive_lcell_comb \ShiftLeft0~31 (
// Equation(s):
// \ShiftLeft0~31_combout  = (Mux301 & (alu_a_mux_output_4)) # (!Mux301 & ((alu_a_mux_output_6)))

	.dataa(gnd),
	.datab(alu_a_mux_output_4),
	.datac(Mux301),
	.datad(alu_a_mux_output_6),
	.cin(gnd),
	.combout(\ShiftLeft0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~31 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N4
cycloneive_lcell_comb \ShiftLeft0~33 (
// Equation(s):
// \ShiftLeft0~33_combout  = (Mux311 & ((\ShiftLeft0~31_combout ))) # (!Mux311 & (\ShiftLeft0~32_combout ))

	.dataa(Mux311),
	.datab(gnd),
	.datac(\ShiftLeft0~32_combout ),
	.datad(\ShiftLeft0~31_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~33 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N14
cycloneive_lcell_comb \ShiftLeft0~30 (
// Equation(s):
// \ShiftLeft0~30_combout  = (\ShiftLeft0~20_combout ) # ((\ShiftLeft0~12_combout  & Mux301))

	.dataa(\ShiftLeft0~12_combout ),
	.datab(gnd),
	.datac(Mux301),
	.datad(\ShiftLeft0~20_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~30 .lut_mask = 16'hFFA0;
defparam \ShiftLeft0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N8
cycloneive_lcell_comb \ShiftLeft0~34 (
// Equation(s):
// \ShiftLeft0~34_combout  = (Mux291 & ((\ShiftLeft0~30_combout ))) # (!Mux291 & (\ShiftLeft0~33_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~33_combout ),
	.datac(Mux291),
	.datad(\ShiftLeft0~30_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~34 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N16
cycloneive_lcell_comb \Mux24~2 (
// Equation(s):
// \Mux24~2_combout  = (!Mux281 & (\Mux19~0_combout  & \ShiftLeft0~34_combout ))

	.dataa(Mux281),
	.datab(gnd),
	.datac(\Mux19~0_combout ),
	.datad(\ShiftLeft0~34_combout ),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~2 .lut_mask = 16'h5000;
defparam \Mux24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N26
cycloneive_lcell_comb \Mux24~3 (
// Equation(s):
// \Mux24~3_combout  = (\Mux27~4_combout  & ((temp_ALUop_output_0 & (\Mux24~1_combout )) # (!temp_ALUop_output_0 & ((\Mux24~2_combout ))))) # (!\Mux27~4_combout  & (((!temp_ALUop_output_0))))

	.dataa(\Mux27~4_combout ),
	.datab(\Mux24~1_combout ),
	.datac(temp_ALUop_output_0),
	.datad(\Mux24~2_combout ),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~3 .lut_mask = 16'h8F85;
defparam \Mux24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N8
cycloneive_lcell_comb \Mux24~4 (
// Equation(s):
// \Mux24~4_combout  = (\Mux24~3_combout  & (((Mux24 & alu_a_mux_output_7)) # (!temp_ALUop_output_1))) # (!\Mux24~3_combout  & (temp_ALUop_output_1 & ((Mux24) # (alu_a_mux_output_7))))

	.dataa(Mux24),
	.datab(alu_a_mux_output_7),
	.datac(\Mux24~3_combout ),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~4 .lut_mask = 16'h8EF0;
defparam \Mux24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N4
cycloneive_lcell_comb \Add0~25 (
// Equation(s):
// \Add0~25_combout  = temp_ALUop_output_0 $ (((temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1) # (temp_imemload_output_7))) # (!temp_ALUsrc_output_0 & (!temp_ALUsrc_output_1))))

	.dataa(temp_ALUsrc_output_0),
	.datab(temp_ALUsrc_output_1),
	.datac(temp_ALUop_output_0),
	.datad(temp_imemload_output_7),
	.cin(gnd),
	.combout(\Add0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~25 .lut_mask = 16'h4B69;
defparam \Add0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N22
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = \Add0~25_combout  $ (((!alu_b_mux_output_7 & (temp_ALUsrc_output_0 $ (!temp_ALUsrc_output_1)))))

	.dataa(temp_ALUsrc_output_0),
	.datab(alu_b_mux_output_7),
	.datac(\Add0~25_combout ),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(\Add0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'hD2E1;
defparam \Add0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N14
cycloneive_lcell_comb \Add0~27 (
// Equation(s):
// \Add0~27_combout  = temp_ALUop_output_0 $ (((temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0))) # (!temp_ALUsrc_output_1 & ((temp_imemload_output_6) # (!temp_ALUsrc_output_0)))))

	.dataa(temp_ALUsrc_output_1),
	.datab(temp_imemload_output_6),
	.datac(temp_ALUop_output_0),
	.datad(temp_ALUsrc_output_0),
	.cin(gnd),
	.combout(\Add0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~27 .lut_mask = 16'h1EA5;
defparam \Add0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N12
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = \Add0~27_combout  $ (((!alu_b_mux_output_6 & (temp_ALUsrc_output_1 $ (!temp_ALUsrc_output_0)))))

	.dataa(temp_ALUsrc_output_1),
	.datab(\Add0~27_combout ),
	.datac(alu_b_mux_output_6),
	.datad(temp_ALUsrc_output_0),
	.cin(gnd),
	.combout(\Add0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'hC6C9;
defparam \Add0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N30
cycloneive_lcell_comb \Add0~29 (
// Equation(s):
// \Add0~29_combout  = (alu_a_mux_output_6 & ((\Add0~28_combout  & (\Add0~24  & VCC)) # (!\Add0~28_combout  & (!\Add0~24 )))) # (!alu_a_mux_output_6 & ((\Add0~28_combout  & (!\Add0~24 )) # (!\Add0~28_combout  & ((\Add0~24 ) # (GND)))))
// \Add0~30  = CARRY((alu_a_mux_output_6 & (!\Add0~28_combout  & !\Add0~24 )) # (!alu_a_mux_output_6 & ((!\Add0~24 ) # (!\Add0~28_combout ))))

	.dataa(alu_a_mux_output_6),
	.datab(\Add0~28_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~24 ),
	.combout(\Add0~29_combout ),
	.cout(\Add0~30 ));
// synopsys translate_off
defparam \Add0~29 .lut_mask = 16'h9617;
defparam \Add0~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N0
cycloneive_lcell_comb \Add0~31 (
// Equation(s):
// \Add0~31_combout  = ((alu_a_mux_output_7 $ (\Add0~26_combout  $ (!\Add0~30 )))) # (GND)
// \Add0~32  = CARRY((alu_a_mux_output_7 & ((\Add0~26_combout ) # (!\Add0~30 ))) # (!alu_a_mux_output_7 & (\Add0~26_combout  & !\Add0~30 )))

	.dataa(alu_a_mux_output_7),
	.datab(\Add0~26_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~30 ),
	.combout(\Add0~31_combout ),
	.cout(\Add0~32 ));
// synopsys translate_off
defparam \Add0~31 .lut_mask = 16'h698E;
defparam \Add0~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N4
cycloneive_lcell_comb \Mux25~5 (
// Equation(s):
// \Mux25~5_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!Mux25 & !alu_a_mux_output_6)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (Mux25 $ (alu_a_mux_output_6))))

	.dataa(Mux25),
	.datab(alu_a_mux_output_6),
	.datac(\Mux19~2_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~5 .lut_mask = 16'hF016;
defparam \Mux25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y43_N30
cycloneive_lcell_comb \ShiftLeft0~18 (
// Equation(s):
// \ShiftLeft0~18_combout  = (!Mux311 & ((Mux301 & (alu_a_mux_output_0)) # (!Mux301 & ((alu_a_mux_output_2)))))

	.dataa(Mux301),
	.datab(Mux311),
	.datac(alu_a_mux_output_0),
	.datad(alu_a_mux_output_2),
	.cin(gnd),
	.combout(\ShiftLeft0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~18 .lut_mask = 16'h3120;
defparam \ShiftLeft0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N6
cycloneive_lcell_comb \ShiftLeft0~104 (
// Equation(s):
// \ShiftLeft0~104_combout  = (\ShiftLeft0~18_combout ) # ((Mux311 & (alu_a_mux_output_1 & !Mux301)))

	.dataa(Mux311),
	.datab(alu_a_mux_output_1),
	.datac(Mux301),
	.datad(\ShiftLeft0~18_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~104 .lut_mask = 16'hFF08;
defparam \ShiftLeft0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N16
cycloneive_lcell_comb \ShiftLeft0~23 (
// Equation(s):
// \ShiftLeft0~23_combout  = (Mux301 & (((alu_a_mux_output_32) # (alu_a_mux_output_3)))) # (!Mux301 & (alu_a_mux_output_5))

	.dataa(Mux301),
	.datab(alu_a_mux_output_5),
	.datac(alu_a_mux_output_32),
	.datad(alu_a_mux_output_3),
	.cin(gnd),
	.combout(\ShiftLeft0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~23 .lut_mask = 16'hEEE4;
defparam \ShiftLeft0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N14
cycloneive_lcell_comb \ShiftLeft0~35 (
// Equation(s):
// \ShiftLeft0~35_combout  = (Mux311 & (\ShiftLeft0~23_combout )) # (!Mux311 & ((\ShiftLeft0~31_combout )))

	.dataa(Mux311),
	.datab(\ShiftLeft0~23_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~31_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~35 .lut_mask = 16'hDD88;
defparam \ShiftLeft0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N28
cycloneive_lcell_comb \ShiftLeft0~36 (
// Equation(s):
// \ShiftLeft0~36_combout  = (Mux291 & (\ShiftLeft0~104_combout )) # (!Mux291 & ((\ShiftLeft0~35_combout )))

	.dataa(Mux291),
	.datab(\ShiftLeft0~104_combout ),
	.datac(\ShiftLeft0~35_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~36 .lut_mask = 16'hD8D8;
defparam \ShiftLeft0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N10
cycloneive_lcell_comb \Mux25~2 (
// Equation(s):
// \Mux25~2_combout  = (!Mux281 & (\Mux19~0_combout  & \ShiftLeft0~36_combout ))

	.dataa(Mux281),
	.datab(gnd),
	.datac(\Mux19~0_combout ),
	.datad(\ShiftLeft0~36_combout ),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~2 .lut_mask = 16'h5000;
defparam \Mux25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N2
cycloneive_lcell_comb \ShiftRight0~61 (
// Equation(s):
// \ShiftRight0~61_combout  = (Mux311 & (\ShiftRight0~60_combout )) # (!Mux311 & ((\ShiftRight0~12_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~60_combout ),
	.datac(Mux311),
	.datad(\ShiftRight0~12_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~61 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N8
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (\Mux27~3_combout  & (\Mux27~2_combout )) # (!\Mux27~3_combout  & ((\Mux27~2_combout  & ((\ShiftRight0~61_combout ))) # (!\Mux27~2_combout  & (\ShiftRight0~58_combout ))))

	.dataa(\Mux27~3_combout ),
	.datab(\Mux27~2_combout ),
	.datac(\ShiftRight0~58_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hDC98;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N16
cycloneive_lcell_comb \ShiftRight0~99 (
// Equation(s):
// \ShiftRight0~99_combout  = (\ShiftRight0~71_combout ) # (\ShiftRight0~72_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftRight0~71_combout ),
	.datad(\ShiftRight0~72_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~99 .lut_mask = 16'hFFF0;
defparam \ShiftRight0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N2
cycloneive_lcell_comb \ShiftRight0~62 (
// Equation(s):
// \ShiftRight0~62_combout  = (!Mux301 & ((Mux311 & ((alu_a_mux_output_15))) # (!Mux311 & (alu_a_mux_output_14))))

	.dataa(Mux311),
	.datab(Mux301),
	.datac(alu_a_mux_output_14),
	.datad(alu_a_mux_output_15),
	.cin(gnd),
	.combout(\ShiftRight0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~62 .lut_mask = 16'h3210;
defparam \ShiftRight0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N30
cycloneive_lcell_comb \ShiftRight0~100 (
// Equation(s):
// \ShiftRight0~100_combout  = (Mux291 & (((\ShiftRight0~99_combout )))) # (!Mux291 & ((\ShiftRight0~63_combout ) # ((\ShiftRight0~62_combout ))))

	.dataa(\ShiftRight0~63_combout ),
	.datab(Mux291),
	.datac(\ShiftRight0~99_combout ),
	.datad(\ShiftRight0~62_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~100 .lut_mask = 16'hF3E2;
defparam \ShiftRight0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N22
cycloneive_lcell_comb \ShiftRight0~101 (
// Equation(s):
// \ShiftRight0~101_combout  = (Mux291 & (((\ShiftRight0~66_combout ) # (\ShiftRight0~65_combout )))) # (!Mux291 & (\ShiftRight0~70_combout ))

	.dataa(\ShiftRight0~70_combout ),
	.datab(\ShiftRight0~66_combout ),
	.datac(Mux291),
	.datad(\ShiftRight0~65_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~101 .lut_mask = 16'hFACA;
defparam \ShiftRight0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N10
cycloneive_lcell_comb \ShiftRight0~102 (
// Equation(s):
// \ShiftRight0~102_combout  = (Mux281 & (\ShiftRight0~44_combout  & (!\ShiftLeft0~13_combout ))) # (!Mux281 & (((\ShiftRight0~101_combout ))))

	.dataa(Mux281),
	.datab(\ShiftRight0~44_combout ),
	.datac(\ShiftLeft0~13_combout ),
	.datad(\ShiftRight0~101_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~102 .lut_mask = 16'h5D08;
defparam \ShiftRight0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N28
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\Mux27~3_combout  & ((\Mux25~0_combout  & ((\ShiftRight0~102_combout ))) # (!\Mux25~0_combout  & (\ShiftRight0~100_combout )))) # (!\Mux27~3_combout  & (\Mux25~0_combout ))

	.dataa(\Mux27~3_combout ),
	.datab(\Mux25~0_combout ),
	.datac(\ShiftRight0~100_combout ),
	.datad(\ShiftRight0~102_combout ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hEC64;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N6
cycloneive_lcell_comb \Mux25~3 (
// Equation(s):
// \Mux25~3_combout  = (temp_ALUop_output_0 & (((\Mux25~1_combout  & \Mux27~4_combout )))) # (!temp_ALUop_output_0 & ((\Mux25~2_combout ) # ((!\Mux27~4_combout ))))

	.dataa(temp_ALUop_output_0),
	.datab(\Mux25~2_combout ),
	.datac(\Mux25~1_combout ),
	.datad(\Mux27~4_combout ),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~3 .lut_mask = 16'hE455;
defparam \Mux25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N6
cycloneive_lcell_comb \Mux25~4 (
// Equation(s):
// \Mux25~4_combout  = (temp_ALUop_output_1 & ((alu_a_mux_output_6 & ((Mux25) # (!\Mux25~3_combout ))) # (!alu_a_mux_output_6 & (!\Mux25~3_combout  & Mux25)))) # (!temp_ALUop_output_1 & (((\Mux25~3_combout ))))

	.dataa(temp_ALUop_output_1),
	.datab(alu_a_mux_output_6),
	.datac(\Mux25~3_combout ),
	.datad(Mux25),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~4 .lut_mask = 16'hDA58;
defparam \Mux25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N14
cycloneive_lcell_comb \ShiftRight0~15 (
// Equation(s):
// \ShiftRight0~15_combout  = (Mux291 & ((\ShiftRight0~11_combout ))) # (!Mux291 & (\ShiftRight0~14_combout ))

	.dataa(gnd),
	.datab(Mux291),
	.datac(\ShiftRight0~14_combout ),
	.datad(\ShiftRight0~11_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~15 .lut_mask = 16'hFC30;
defparam \ShiftRight0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N28
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = ((\ShiftLeft0~10_combout ) # ((\ShiftLeft0~26_combout ) # (Mux271))) # (!temp_ALUop_output_0)

	.dataa(temp_ALUop_output_0),
	.datab(\ShiftLeft0~10_combout ),
	.datac(\ShiftLeft0~26_combout ),
	.datad(Mux271),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'hFFFD;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N24
cycloneive_lcell_comb \ShiftRight0~25 (
// Equation(s):
// \ShiftRight0~25_combout  = (Mux301 & ((Mux311 & ((alu_a_mux_output_24))) # (!Mux311 & (alu_a_mux_output_23))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_23),
	.datac(alu_a_mux_output_24),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftRight0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~25 .lut_mask = 16'hA088;
defparam \ShiftRight0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N26
cycloneive_lcell_comb \ShiftRight0~27 (
// Equation(s):
// \ShiftRight0~27_combout  = (Mux291 & ((\ShiftRight0~26_combout ) # ((\ShiftRight0~25_combout )))) # (!Mux291 & (((\ShiftRight0~24_combout ))))

	.dataa(Mux291),
	.datab(\ShiftRight0~26_combout ),
	.datac(\ShiftRight0~25_combout ),
	.datad(\ShiftRight0~24_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~27 .lut_mask = 16'hFDA8;
defparam \ShiftRight0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N30
cycloneive_lcell_comb \ShiftLeft0~37 (
// Equation(s):
// \ShiftLeft0~37_combout  = (Mux301 & ((alu_a_mux_output_6))) # (!Mux301 & (alu_a_mux_output_8))

	.dataa(gnd),
	.datab(Mux301),
	.datac(alu_a_mux_output_8),
	.datad(alu_a_mux_output_6),
	.cin(gnd),
	.combout(\ShiftLeft0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~37 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N8
cycloneive_lcell_comb \ShiftLeft0~39 (
// Equation(s):
// \ShiftLeft0~39_combout  = (Mux311 & ((\ShiftLeft0~37_combout ))) # (!Mux311 & (\ShiftLeft0~38_combout ))

	.dataa(\ShiftLeft0~38_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~37_combout ),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftLeft0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~39 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N16
cycloneive_lcell_comb \ShiftLeft0~24 (
// Equation(s):
// \ShiftLeft0~24_combout  = (Mux311 & ((\ShiftLeft0~22_combout ))) # (!Mux311 & (\ShiftLeft0~23_combout ))

	.dataa(Mux311),
	.datab(\ShiftLeft0~23_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~22_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~24 .lut_mask = 16'hEE44;
defparam \ShiftLeft0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N6
cycloneive_lcell_comb \ShiftLeft0~40 (
// Equation(s):
// \ShiftLeft0~40_combout  = (Mux291 & ((\ShiftLeft0~24_combout ))) # (!Mux291 & (\ShiftLeft0~39_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~39_combout ),
	.datac(Mux291),
	.datad(\ShiftLeft0~24_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~40 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N6
cycloneive_lcell_comb \ShiftLeft0~41 (
// Equation(s):
// \ShiftLeft0~41_combout  = (Mux281 & (!\ShiftLeft0~13_combout  & (\ShiftLeft0~12_combout ))) # (!Mux281 & (((\ShiftLeft0~40_combout ))))

	.dataa(\ShiftLeft0~13_combout ),
	.datab(\ShiftLeft0~12_combout ),
	.datac(\ShiftLeft0~40_combout ),
	.datad(Mux281),
	.cin(gnd),
	.combout(\ShiftLeft0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~41 .lut_mask = 16'h44F0;
defparam \ShiftLeft0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N24
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (!\ShiftLeft0~26_combout  & (!\ShiftLeft0~10_combout  & (!Mux271 & \ShiftLeft0~41_combout )))

	.dataa(\ShiftLeft0~26_combout ),
	.datab(\ShiftLeft0~10_combout ),
	.datac(Mux271),
	.datad(\ShiftLeft0~41_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'h0100;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N28
cycloneive_lcell_comb \Mux19~4 (
// Equation(s):
// \Mux19~4_combout  = ((!\Mux19~0_combout  & !\ShiftLeft0~11_combout )) # (!temp_ALUop_output_0)

	.dataa(gnd),
	.datab(\Mux19~0_combout ),
	.datac(temp_ALUop_output_0),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\Mux19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~4 .lut_mask = 16'h0F3F;
defparam \Mux19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N0
cycloneive_lcell_comb \Mux19~5 (
// Equation(s):
// \Mux19~5_combout  = (temp_ALUop_output_0 & ((Mux281) # (!\Mux19~0_combout )))

	.dataa(temp_ALUop_output_0),
	.datab(gnd),
	.datac(\Mux19~0_combout ),
	.datad(Mux281),
	.cin(gnd),
	.combout(\Mux19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~5 .lut_mask = 16'hAA0A;
defparam \Mux19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N12
cycloneive_lcell_comb \Mux22~2 (
// Equation(s):
// \Mux22~2_combout  = (\Mux19~4_combout  & ((\Mux19~5_combout  & (\ShiftRight0~103_combout )) # (!\Mux19~5_combout  & ((\Mux22~1_combout ))))) # (!\Mux19~4_combout  & (((!\Mux19~5_combout ))))

	.dataa(\ShiftRight0~103_combout ),
	.datab(\Mux22~1_combout ),
	.datac(\Mux19~4_combout ),
	.datad(\Mux19~5_combout ),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~2 .lut_mask = 16'hA0CF;
defparam \Mux22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N14
cycloneive_lcell_comb \Mux22~3 (
// Equation(s):
// \Mux22~3_combout  = (\Mux19~3_combout  & (((\Mux22~2_combout )))) # (!\Mux19~3_combout  & ((\Mux22~2_combout  & (\ShiftRight0~15_combout )) # (!\Mux22~2_combout  & ((\ShiftRight0~27_combout )))))

	.dataa(\ShiftRight0~15_combout ),
	.datab(\Mux19~3_combout ),
	.datac(\ShiftRight0~27_combout ),
	.datad(\Mux22~2_combout ),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~3 .lut_mask = 16'hEE30;
defparam \Mux22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N6
cycloneive_lcell_comb \Add0~33 (
// Equation(s):
// \Add0~33_combout  = temp_ALUop_output_0 $ (Mux22)

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(Mux22),
	.cin(gnd),
	.combout(\Add0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~33 .lut_mask = 16'h0FF0;
defparam \Add0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N28
cycloneive_lcell_comb \Add0~34 (
// Equation(s):
// \Add0~34_combout  = temp_ALUop_output_0 $ (Mux23)

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(Mux23),
	.cin(gnd),
	.combout(\Add0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~34 .lut_mask = 16'h0FF0;
defparam \Add0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N2
cycloneive_lcell_comb \Add0~35 (
// Equation(s):
// \Add0~35_combout  = (alu_a_mux_output_8 & ((\Add0~34_combout  & (\Add0~32  & VCC)) # (!\Add0~34_combout  & (!\Add0~32 )))) # (!alu_a_mux_output_8 & ((\Add0~34_combout  & (!\Add0~32 )) # (!\Add0~34_combout  & ((\Add0~32 ) # (GND)))))
// \Add0~36  = CARRY((alu_a_mux_output_8 & (!\Add0~34_combout  & !\Add0~32 )) # (!alu_a_mux_output_8 & ((!\Add0~32 ) # (!\Add0~34_combout ))))

	.dataa(alu_a_mux_output_8),
	.datab(\Add0~34_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~32 ),
	.combout(\Add0~35_combout ),
	.cout(\Add0~36 ));
// synopsys translate_off
defparam \Add0~35 .lut_mask = 16'h9617;
defparam \Add0~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N4
cycloneive_lcell_comb \Add0~37 (
// Equation(s):
// \Add0~37_combout  = ((\Add0~33_combout  $ (alu_a_mux_output_9 $ (!\Add0~36 )))) # (GND)
// \Add0~38  = CARRY((\Add0~33_combout  & ((alu_a_mux_output_9) # (!\Add0~36 ))) # (!\Add0~33_combout  & (alu_a_mux_output_9 & !\Add0~36 )))

	.dataa(\Add0~33_combout ),
	.datab(alu_a_mux_output_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~36 ),
	.combout(\Add0~37_combout ),
	.cout(\Add0~38 ));
// synopsys translate_off
defparam \Add0~37 .lut_mask = 16'h698E;
defparam \Add0~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N12
cycloneive_lcell_comb \Mux22~4 (
// Equation(s):
// \Mux22~4_combout  = (\Mux19~1_combout  & (((\Mux19~2_combout )))) # (!\Mux19~1_combout  & ((Mux22 & (!alu_a_mux_output_9 & !\Mux19~2_combout )) # (!Mux22 & (alu_a_mux_output_9 $ (\Mux19~2_combout )))))

	.dataa(\Mux19~1_combout ),
	.datab(Mux22),
	.datac(alu_a_mux_output_9),
	.datad(\Mux19~2_combout ),
	.cin(gnd),
	.combout(\Mux22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~4 .lut_mask = 16'hAB14;
defparam \Mux22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N26
cycloneive_lcell_comb \Mux23~4 (
// Equation(s):
// \Mux23~4_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!alu_a_mux_output_8 & !Mux23)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (alu_a_mux_output_8 $ (Mux23))))

	.dataa(alu_a_mux_output_8),
	.datab(\Mux19~2_combout ),
	.datac(Mux23),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~4 .lut_mask = 16'hCC16;
defparam \Mux23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N16
cycloneive_lcell_comb \ShiftRight0~38 (
// Equation(s):
// \ShiftRight0~38_combout  = (Mux311 & (\ShiftRight0~10_combout )) # (!Mux311 & ((\ShiftRight0~37_combout )))

	.dataa(gnd),
	.datab(Mux311),
	.datac(\ShiftRight0~10_combout ),
	.datad(\ShiftRight0~37_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~38 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N6
cycloneive_lcell_comb \ShiftRight0~41 (
// Equation(s):
// \ShiftRight0~41_combout  = (Mux291 & (\ShiftRight0~38_combout )) # (!Mux291 & ((\ShiftRight0~40_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~38_combout ),
	.datac(Mux291),
	.datad(\ShiftRight0~40_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~41 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N22
cycloneive_lcell_comb \ShiftRight0~47 (
// Equation(s):
// \ShiftRight0~47_combout  = (Mux301 & ((Mux311 & ((alu_a_mux_output_23))) # (!Mux311 & (alu_a_mux_output_22))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_22),
	.datac(alu_a_mux_output_23),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftRight0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~47 .lut_mask = 16'hA088;
defparam \ShiftRight0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N4
cycloneive_lcell_comb \ShiftRight0~48 (
// Equation(s):
// \ShiftRight0~48_combout  = (\ShiftRight0~47_combout ) # (\ShiftRight0~46_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftRight0~47_combout ),
	.datad(\ShiftRight0~46_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~48 .lut_mask = 16'hFFF0;
defparam \ShiftRight0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N2
cycloneive_lcell_comb \ShiftRight0~49 (
// Equation(s):
// \ShiftRight0~49_combout  = (!Mux301 & ((Mux311 & ((alu_a_mux_output_17))) # (!Mux311 & (alu_a_mux_output_16))))

	.dataa(Mux311),
	.datab(alu_a_mux_output_16),
	.datac(Mux301),
	.datad(alu_a_mux_output_17),
	.cin(gnd),
	.combout(\ShiftRight0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~49 .lut_mask = 16'h0E04;
defparam \ShiftRight0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N26
cycloneive_lcell_comb \ShiftRight0~51 (
// Equation(s):
// \ShiftRight0~51_combout  = (Mux291 & (((\ShiftRight0~48_combout )))) # (!Mux291 & ((\ShiftRight0~50_combout ) # ((\ShiftRight0~49_combout ))))

	.dataa(\ShiftRight0~50_combout ),
	.datab(\ShiftRight0~48_combout ),
	.datac(Mux291),
	.datad(\ShiftRight0~49_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~51 .lut_mask = 16'hCFCA;
defparam \ShiftRight0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y40_N24
cycloneive_lcell_comb \ShiftLeft0~43 (
// Equation(s):
// \ShiftLeft0~43_combout  = (!Mux311 & ((Mux301 & ((alu_a_mux_output_6))) # (!Mux301 & (alu_a_mux_output_8))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_8),
	.datac(alu_a_mux_output_6),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftLeft0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~43 .lut_mask = 16'h00E4;
defparam \ShiftLeft0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N22
cycloneive_lcell_comb \ShiftLeft0~44 (
// Equation(s):
// \ShiftLeft0~44_combout  = (Mux291 & (((\ShiftLeft0~28_combout )))) # (!Mux291 & ((\ShiftLeft0~42_combout ) # ((\ShiftLeft0~43_combout ))))

	.dataa(\ShiftLeft0~42_combout ),
	.datab(\ShiftLeft0~28_combout ),
	.datac(Mux291),
	.datad(\ShiftLeft0~43_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~44 .lut_mask = 16'hCFCA;
defparam \ShiftLeft0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N0
cycloneive_lcell_comb \ShiftLeft0~45 (
// Equation(s):
// \ShiftLeft0~45_combout  = (Mux281 & (!Mux291 & ((\ShiftLeft0~16_combout )))) # (!Mux281 & (((\ShiftLeft0~44_combout ))))

	.dataa(Mux291),
	.datab(Mux281),
	.datac(\ShiftLeft0~44_combout ),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~45 .lut_mask = 16'h7430;
defparam \ShiftLeft0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N2
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (!Mux271 & (!\ShiftLeft0~26_combout  & (!\ShiftLeft0~10_combout  & \ShiftLeft0~45_combout )))

	.dataa(Mux271),
	.datab(\ShiftLeft0~26_combout ),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\ShiftLeft0~45_combout ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'h0100;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N0
cycloneive_lcell_comb \Mux23~2 (
// Equation(s):
// \Mux23~2_combout  = (\Mux19~4_combout  & ((\Mux19~5_combout  & (\ShiftRight0~104_combout )) # (!\Mux19~5_combout  & ((\Mux23~1_combout ))))) # (!\Mux19~4_combout  & (((!\Mux19~5_combout ))))

	.dataa(\ShiftRight0~104_combout ),
	.datab(\Mux23~1_combout ),
	.datac(\Mux19~4_combout ),
	.datad(\Mux19~5_combout ),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~2 .lut_mask = 16'hA0CF;
defparam \Mux23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N24
cycloneive_lcell_comb \Mux23~3 (
// Equation(s):
// \Mux23~3_combout  = (\Mux19~3_combout  & (((\Mux23~2_combout )))) # (!\Mux19~3_combout  & ((\Mux23~2_combout  & (\ShiftRight0~41_combout )) # (!\Mux23~2_combout  & ((\ShiftRight0~51_combout )))))

	.dataa(\ShiftRight0~41_combout ),
	.datab(\Mux19~3_combout ),
	.datac(\ShiftRight0~51_combout ),
	.datad(\Mux23~2_combout ),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~3 .lut_mask = 16'hEE30;
defparam \Mux23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y43_N12
cycloneive_lcell_comb \Mux20~4 (
// Equation(s):
// \Mux20~4_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!alu_a_mux_output_11 & !Mux20)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (alu_a_mux_output_11 $ (Mux20))))

	.dataa(alu_a_mux_output_11),
	.datab(\Mux19~2_combout ),
	.datac(\Mux19~1_combout ),
	.datad(Mux20),
	.cin(gnd),
	.combout(\Mux20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~4 .lut_mask = 16'hC1C6;
defparam \Mux20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N22
cycloneive_lcell_comb \Add0~39 (
// Equation(s):
// \Add0~39_combout  = temp_ALUop_output_0 $ (Mux20)

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(Mux20),
	.cin(gnd),
	.combout(\Add0~39_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~39 .lut_mask = 16'h0FF0;
defparam \Add0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N24
cycloneive_lcell_comb \Add0~40 (
// Equation(s):
// \Add0~40_combout  = temp_ALUop_output_0 $ (Mux21)

	.dataa(gnd),
	.datab(temp_ALUop_output_0),
	.datac(gnd),
	.datad(Mux21),
	.cin(gnd),
	.combout(\Add0~40_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~40 .lut_mask = 16'h33CC;
defparam \Add0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N6
cycloneive_lcell_comb \Add0~41 (
// Equation(s):
// \Add0~41_combout  = (alu_a_mux_output_10 & ((\Add0~40_combout  & (\Add0~38  & VCC)) # (!\Add0~40_combout  & (!\Add0~38 )))) # (!alu_a_mux_output_10 & ((\Add0~40_combout  & (!\Add0~38 )) # (!\Add0~40_combout  & ((\Add0~38 ) # (GND)))))
// \Add0~42  = CARRY((alu_a_mux_output_10 & (!\Add0~40_combout  & !\Add0~38 )) # (!alu_a_mux_output_10 & ((!\Add0~38 ) # (!\Add0~40_combout ))))

	.dataa(alu_a_mux_output_10),
	.datab(\Add0~40_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~38 ),
	.combout(\Add0~41_combout ),
	.cout(\Add0~42 ));
// synopsys translate_off
defparam \Add0~41 .lut_mask = 16'h9617;
defparam \Add0~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N8
cycloneive_lcell_comb \Add0~43 (
// Equation(s):
// \Add0~43_combout  = ((\Add0~39_combout  $ (alu_a_mux_output_11 $ (!\Add0~42 )))) # (GND)
// \Add0~44  = CARRY((\Add0~39_combout  & ((alu_a_mux_output_11) # (!\Add0~42 ))) # (!\Add0~39_combout  & (alu_a_mux_output_11 & !\Add0~42 )))

	.dataa(\Add0~39_combout ),
	.datab(alu_a_mux_output_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~42 ),
	.combout(\Add0~43_combout ),
	.cout(\Add0~44 ));
// synopsys translate_off
defparam \Add0~43 .lut_mask = 16'h698E;
defparam \Add0~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N16
cycloneive_lcell_comb \ShiftRight0~83 (
// Equation(s):
// \ShiftRight0~83_combout  = (Mux291 & (\ShiftRight0~80_combout )) # (!Mux291 & (((\ShiftRight0~81_combout ) # (\ShiftRight0~82_combout ))))

	.dataa(Mux291),
	.datab(\ShiftRight0~80_combout ),
	.datac(\ShiftRight0~81_combout ),
	.datad(\ShiftRight0~82_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~83 .lut_mask = 16'hDDD8;
defparam \ShiftRight0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N0
cycloneive_lcell_comb \ShiftRight0~105 (
// Equation(s):
// \ShiftRight0~105_combout  = (!Mux281 & \ShiftRight0~83_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux281),
	.datad(\ShiftRight0~83_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~105_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~105 .lut_mask = 16'h0F00;
defparam \ShiftRight0~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N26
cycloneive_lcell_comb \Mux20~2 (
// Equation(s):
// \Mux20~2_combout  = (\Mux19~4_combout  & ((\Mux19~5_combout  & ((\ShiftRight0~105_combout ))) # (!\Mux19~5_combout  & (\Mux20~1_combout )))) # (!\Mux19~4_combout  & (((!\Mux19~5_combout ))))

	.dataa(\Mux20~1_combout ),
	.datab(\Mux19~4_combout ),
	.datac(\Mux19~5_combout ),
	.datad(\ShiftRight0~105_combout ),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~2 .lut_mask = 16'hCB0B;
defparam \Mux20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N28
cycloneive_lcell_comb \ShiftRight0~84 (
// Equation(s):
// \ShiftRight0~84_combout  = (Mux311 & ((alu_a_mux_output_26) # ((!Mux301)))) # (!Mux311 & (((Mux301 & alu_a_mux_output_25))))

	.dataa(Mux311),
	.datab(alu_a_mux_output_26),
	.datac(Mux301),
	.datad(alu_a_mux_output_25),
	.cin(gnd),
	.combout(\ShiftRight0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~84 .lut_mask = 16'hDA8A;
defparam \ShiftRight0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N26
cycloneive_lcell_comb \ShiftRight0~85 (
// Equation(s):
// \ShiftRight0~85_combout  = (Mux301 & (((\ShiftRight0~84_combout )))) # (!Mux301 & ((\ShiftRight0~84_combout  & ((alu_a_mux_output_24))) # (!\ShiftRight0~84_combout  & (alu_a_mux_output_23))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_23),
	.datac(alu_a_mux_output_24),
	.datad(\ShiftRight0~84_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~85 .lut_mask = 16'hFA44;
defparam \ShiftRight0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N20
cycloneive_lcell_comb \ShiftRight0~86 (
// Equation(s):
// \ShiftRight0~86_combout  = (Mux301 & ((Mux311 & ((alu_a_mux_output_22))) # (!Mux311 & (alu_a_mux_output_21)))) # (!Mux301 & (((Mux311))))

	.dataa(alu_a_mux_output_21),
	.datab(Mux301),
	.datac(Mux311),
	.datad(alu_a_mux_output_22),
	.cin(gnd),
	.combout(\ShiftRight0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~86 .lut_mask = 16'hF838;
defparam \ShiftRight0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N18
cycloneive_lcell_comb \ShiftRight0~87 (
// Equation(s):
// \ShiftRight0~87_combout  = (Mux301 & (((\ShiftRight0~86_combout )))) # (!Mux301 & ((\ShiftRight0~86_combout  & (alu_a_mux_output_20)) # (!\ShiftRight0~86_combout  & ((alu_a_mux_output_19)))))

	.dataa(alu_a_mux_output_20),
	.datab(Mux301),
	.datac(alu_a_mux_output_19),
	.datad(\ShiftRight0~86_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~87 .lut_mask = 16'hEE30;
defparam \ShiftRight0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N30
cycloneive_lcell_comb \ShiftRight0~88 (
// Equation(s):
// \ShiftRight0~88_combout  = (Mux291 & (\ShiftRight0~85_combout )) # (!Mux291 & ((\ShiftRight0~87_combout )))

	.dataa(Mux291),
	.datab(gnd),
	.datac(\ShiftRight0~85_combout ),
	.datad(\ShiftRight0~87_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~88 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N28
cycloneive_lcell_comb \Mux20~3 (
// Equation(s):
// \Mux20~3_combout  = (\Mux20~2_combout  & ((\ShiftRight0~79_combout ) # ((\Mux19~3_combout )))) # (!\Mux20~2_combout  & (((\ShiftRight0~88_combout  & !\Mux19~3_combout ))))

	.dataa(\Mux20~2_combout ),
	.datab(\ShiftRight0~79_combout ),
	.datac(\ShiftRight0~88_combout ),
	.datad(\Mux19~3_combout ),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~3 .lut_mask = 16'hAAD8;
defparam \Mux20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N26
cycloneive_lcell_comb \ShiftRight0~64 (
// Equation(s):
// \ShiftRight0~64_combout  = (Mux291 & ((\ShiftRight0~63_combout ) # ((\ShiftRight0~62_combout )))) # (!Mux291 & (((\ShiftRight0~61_combout ))))

	.dataa(\ShiftRight0~63_combout ),
	.datab(\ShiftRight0~61_combout ),
	.datac(Mux291),
	.datad(\ShiftRight0~62_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~64 .lut_mask = 16'hFCAC;
defparam \ShiftRight0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N8
cycloneive_lcell_comb \ShiftLeft0~46 (
// Equation(s):
// \ShiftLeft0~46_combout  = (Mux301 & (alu_a_mux_output_8)) # (!Mux301 & ((alu_a_mux_output_10)))

	.dataa(alu_a_mux_output_8),
	.datab(gnd),
	.datac(alu_a_mux_output_10),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftLeft0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~46 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N4
cycloneive_lcell_comb \ShiftLeft0~51 (
// Equation(s):
// \ShiftLeft0~51_combout  = (Mux311 & (\ShiftLeft0~38_combout )) # (!Mux311 & ((\ShiftLeft0~46_combout )))

	.dataa(\ShiftLeft0~38_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~46_combout ),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftLeft0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~51 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N10
cycloneive_lcell_comb \ShiftLeft0~52 (
// Equation(s):
// \ShiftLeft0~52_combout  = (Mux291 & (\ShiftLeft0~35_combout )) # (!Mux291 & ((\ShiftLeft0~51_combout )))

	.dataa(Mux291),
	.datab(\ShiftLeft0~35_combout ),
	.datac(\ShiftLeft0~51_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~52 .lut_mask = 16'hD8D8;
defparam \ShiftLeft0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N20
cycloneive_lcell_comb \ShiftLeft0~53 (
// Equation(s):
// \ShiftLeft0~53_combout  = (Mux281 & (!Mux291 & (\ShiftLeft0~104_combout ))) # (!Mux281 & (((\ShiftLeft0~52_combout ))))

	.dataa(Mux291),
	.datab(\ShiftLeft0~104_combout ),
	.datac(Mux281),
	.datad(\ShiftLeft0~52_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~53 .lut_mask = 16'h4F40;
defparam \ShiftLeft0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N12
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (!\ShiftLeft0~26_combout  & (!\ShiftLeft0~10_combout  & (!Mux271 & \ShiftLeft0~53_combout )))

	.dataa(\ShiftLeft0~26_combout ),
	.datab(\ShiftLeft0~10_combout ),
	.datac(Mux271),
	.datad(\ShiftLeft0~53_combout ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'h0100;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N22
cycloneive_lcell_comb \Mux21~2 (
// Equation(s):
// \Mux21~2_combout  = (\Mux19~4_combout  & ((\Mux19~5_combout  & (\ShiftRight0~107_combout )) # (!\Mux19~5_combout  & ((\Mux21~1_combout ))))) # (!\Mux19~4_combout  & (((!\Mux19~5_combout ))))

	.dataa(\ShiftRight0~107_combout ),
	.datab(\Mux21~1_combout ),
	.datac(\Mux19~4_combout ),
	.datad(\Mux19~5_combout ),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~2 .lut_mask = 16'hA0CF;
defparam \Mux21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N4
cycloneive_lcell_comb \Mux21~3 (
// Equation(s):
// \Mux21~3_combout  = (\Mux19~3_combout  & (((\Mux21~2_combout )))) # (!\Mux19~3_combout  & ((\Mux21~2_combout  & ((\ShiftRight0~64_combout ))) # (!\Mux21~2_combout  & (\ShiftRight0~73_combout ))))

	.dataa(\ShiftRight0~73_combout ),
	.datab(\Mux19~3_combout ),
	.datac(\ShiftRight0~64_combout ),
	.datad(\Mux21~2_combout ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~3 .lut_mask = 16'hFC22;
defparam \Mux21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y43_N0
cycloneive_lcell_comb \Mux21~4 (
// Equation(s):
// \Mux21~4_combout  = (\Mux19~1_combout  & (((\Mux19~2_combout )))) # (!\Mux19~1_combout  & ((Mux21 & (!\Mux19~2_combout  & !alu_a_mux_output_10)) # (!Mux21 & (\Mux19~2_combout  $ (alu_a_mux_output_10)))))

	.dataa(Mux21),
	.datab(\Mux19~1_combout ),
	.datac(\Mux19~2_combout ),
	.datad(alu_a_mux_output_10),
	.cin(gnd),
	.combout(\Mux21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~4 .lut_mask = 16'hC1D2;
defparam \Mux21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N18
cycloneive_lcell_comb \Add0~45 (
// Equation(s):
// \Add0~45_combout  = temp_ALUop_output_0 $ (Mux18)

	.dataa(temp_ALUop_output_0),
	.datab(Mux18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add0~45_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~45 .lut_mask = 16'h6666;
defparam \Add0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N10
cycloneive_lcell_comb \Add0~47 (
// Equation(s):
// \Add0~47_combout  = (\Add0~46_combout  & ((alu_a_mux_output_12 & (\Add0~44  & VCC)) # (!alu_a_mux_output_12 & (!\Add0~44 )))) # (!\Add0~46_combout  & ((alu_a_mux_output_12 & (!\Add0~44 )) # (!alu_a_mux_output_12 & ((\Add0~44 ) # (GND)))))
// \Add0~48  = CARRY((\Add0~46_combout  & (!alu_a_mux_output_12 & !\Add0~44 )) # (!\Add0~46_combout  & ((!\Add0~44 ) # (!alu_a_mux_output_12))))

	.dataa(\Add0~46_combout ),
	.datab(alu_a_mux_output_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~44 ),
	.combout(\Add0~47_combout ),
	.cout(\Add0~48 ));
// synopsys translate_off
defparam \Add0~47 .lut_mask = 16'h9617;
defparam \Add0~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N12
cycloneive_lcell_comb \Add0~49 (
// Equation(s):
// \Add0~49_combout  = ((\Add0~45_combout  $ (alu_a_mux_output_13 $ (!\Add0~48 )))) # (GND)
// \Add0~50  = CARRY((\Add0~45_combout  & ((alu_a_mux_output_13) # (!\Add0~48 ))) # (!\Add0~45_combout  & (alu_a_mux_output_13 & !\Add0~48 )))

	.dataa(\Add0~45_combout ),
	.datab(alu_a_mux_output_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~48 ),
	.combout(\Add0~49_combout ),
	.cout(\Add0~50 ));
// synopsys translate_off
defparam \Add0~49 .lut_mask = 16'h698E;
defparam \Add0~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N8
cycloneive_lcell_comb \ShiftLeft0~55 (
// Equation(s):
// \ShiftLeft0~55_combout  = (Mux301 & ((alu_a_mux_output_11))) # (!Mux301 & (alu_a_mux_output_13))

	.dataa(alu_a_mux_output_13),
	.datab(gnd),
	.datac(alu_a_mux_output_11),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftLeft0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~55 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N10
cycloneive_lcell_comb \ShiftLeft0~54 (
// Equation(s):
// \ShiftLeft0~54_combout  = (Mux301 & (alu_a_mux_output_10)) # (!Mux301 & ((alu_a_mux_output_12)))

	.dataa(Mux301),
	.datab(gnd),
	.datac(alu_a_mux_output_10),
	.datad(alu_a_mux_output_12),
	.cin(gnd),
	.combout(\ShiftLeft0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~54 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N22
cycloneive_lcell_comb \ShiftLeft0~56 (
// Equation(s):
// \ShiftLeft0~56_combout  = (Mux311 & ((\ShiftLeft0~54_combout ))) # (!Mux311 & (\ShiftLeft0~55_combout ))

	.dataa(gnd),
	.datab(Mux311),
	.datac(\ShiftLeft0~55_combout ),
	.datad(\ShiftLeft0~54_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~56 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N30
cycloneive_lcell_comb \ShiftLeft0~57 (
// Equation(s):
// \ShiftLeft0~57_combout  = (Mux291 & (\ShiftLeft0~39_combout )) # (!Mux291 & ((\ShiftLeft0~56_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~39_combout ),
	.datac(Mux291),
	.datad(\ShiftLeft0~56_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~57 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N2
cycloneive_lcell_comb \ShiftLeft0~25 (
// Equation(s):
// \ShiftLeft0~25_combout  = (Mux291 & (!Mux301 & (\ShiftLeft0~12_combout ))) # (!Mux291 & (((\ShiftLeft0~24_combout ))))

	.dataa(Mux301),
	.datab(\ShiftLeft0~12_combout ),
	.datac(Mux291),
	.datad(\ShiftLeft0~24_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~25 .lut_mask = 16'h4F40;
defparam \ShiftLeft0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N14
cycloneive_lcell_comb \ShiftLeft0~58 (
// Equation(s):
// \ShiftLeft0~58_combout  = (Mux281 & ((\ShiftLeft0~25_combout ))) # (!Mux281 & (\ShiftLeft0~57_combout ))

	.dataa(Mux281),
	.datab(gnd),
	.datac(\ShiftLeft0~57_combout ),
	.datad(\ShiftLeft0~25_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~58 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N14
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (!\ShiftLeft0~26_combout  & (!Mux271 & (!\ShiftLeft0~10_combout  & \ShiftLeft0~58_combout )))

	.dataa(\ShiftLeft0~26_combout ),
	.datab(Mux271),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\ShiftLeft0~58_combout ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'h0100;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N28
cycloneive_lcell_comb \ShiftRight0~17 (
// Equation(s):
// \ShiftRight0~17_combout  = (Mux301 & (((alu_a_mux_output_311 & !Mux311)))) # (!Mux301 & (alu_a_mux_output_30 & ((Mux311))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_30),
	.datac(alu_a_mux_output_311),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftRight0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~17 .lut_mask = 16'h44A0;
defparam \ShiftRight0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N26
cycloneive_lcell_comb \ShiftRight0~18 (
// Equation(s):
// \ShiftRight0~18_combout  = (\ShiftRight0~17_combout ) # ((!Mux311 & (alu_a_mux_output_29 & !Mux301)))

	.dataa(Mux311),
	.datab(\ShiftRight0~17_combout ),
	.datac(alu_a_mux_output_29),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftRight0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~18 .lut_mask = 16'hCCDC;
defparam \ShiftRight0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N0
cycloneive_lcell_comb \ShiftRight0~111 (
// Equation(s):
// \ShiftRight0~111_combout  = (!Mux281 & (!Mux291 & \ShiftRight0~18_combout ))

	.dataa(gnd),
	.datab(Mux281),
	.datac(Mux291),
	.datad(\ShiftRight0~18_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~111_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~111 .lut_mask = 16'h0300;
defparam \ShiftRight0~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N8
cycloneive_lcell_comb \Mux18~2 (
// Equation(s):
// \Mux18~2_combout  = (\Mux19~5_combout  & (((\Mux19~4_combout  & \ShiftRight0~111_combout )))) # (!\Mux19~5_combout  & ((\Mux18~1_combout ) # ((!\Mux19~4_combout ))))

	.dataa(\Mux19~5_combout ),
	.datab(\Mux18~1_combout ),
	.datac(\Mux19~4_combout ),
	.datad(\ShiftRight0~111_combout ),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~2 .lut_mask = 16'hE545;
defparam \Mux18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N10
cycloneive_lcell_comb \Mux18~3 (
// Equation(s):
// \Mux18~3_combout  = (\Mux19~3_combout  & (((\Mux18~2_combout )))) # (!\Mux19~3_combout  & ((\Mux18~2_combout  & ((\ShiftRight0~90_combout ))) # (!\Mux18~2_combout  & (\ShiftRight0~91_combout ))))

	.dataa(\Mux19~3_combout ),
	.datab(\ShiftRight0~91_combout ),
	.datac(\Mux18~2_combout ),
	.datad(\ShiftRight0~90_combout ),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~3 .lut_mask = 16'hF4A4;
defparam \Mux18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N2
cycloneive_lcell_comb \Mux18~4 (
// Equation(s):
// \Mux18~4_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!Mux18 & !alu_a_mux_output_13)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (Mux18 $ (alu_a_mux_output_13))))

	.dataa(Mux18),
	.datab(alu_a_mux_output_13),
	.datac(\Mux19~2_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~4 .lut_mask = 16'hF016;
defparam \Mux18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N4
cycloneive_lcell_comb \Add0~46 (
// Equation(s):
// \Add0~46_combout  = temp_ALUop_output_0 $ (Mux19)

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(Mux19),
	.cin(gnd),
	.combout(\Add0~46_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~46 .lut_mask = 16'h0FF0;
defparam \Add0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N28
cycloneive_lcell_comb \Mux19~11 (
// Equation(s):
// \Mux19~11_combout  = (\Mux19~1_combout  & (((\Mux19~2_combout )))) # (!\Mux19~1_combout  & ((alu_a_mux_output_12 & (!\Mux19~2_combout  & !Mux19)) # (!alu_a_mux_output_12 & (\Mux19~2_combout  $ (Mux19)))))

	.dataa(alu_a_mux_output_12),
	.datab(\Mux19~1_combout ),
	.datac(\Mux19~2_combout ),
	.datad(Mux19),
	.cin(gnd),
	.combout(\Mux19~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~11 .lut_mask = 16'hC1D2;
defparam \Mux19~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N6
cycloneive_lcell_comb \ShiftRight0~93 (
// Equation(s):
// \ShiftRight0~93_combout  = (Mux291 & ((\ShiftRight0~50_combout ) # ((\ShiftRight0~49_combout )))) # (!Mux291 & (((\ShiftRight0~38_combout ))))

	.dataa(\ShiftRight0~50_combout ),
	.datab(\ShiftRight0~38_combout ),
	.datac(Mux291),
	.datad(\ShiftRight0~49_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~93 .lut_mask = 16'hFCAC;
defparam \ShiftRight0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N22
cycloneive_lcell_comb \ShiftRight0~108 (
// Equation(s):
// \ShiftRight0~108_combout  = (\ShiftRight0~59_combout  & ((\ShiftRight0~43_combout ) # ((Mux301 & \ShiftRight0~44_combout ))))

	.dataa(\ShiftRight0~59_combout ),
	.datab(\ShiftRight0~43_combout ),
	.datac(Mux301),
	.datad(\ShiftRight0~44_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~108_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~108 .lut_mask = 16'hA888;
defparam \ShiftRight0~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N30
cycloneive_lcell_comb \Mux19~9 (
// Equation(s):
// \Mux19~9_combout  = (\Mux19~4_combout  & ((\Mux19~5_combout  & ((\ShiftRight0~108_combout ))) # (!\Mux19~5_combout  & (\Mux19~8_combout )))) # (!\Mux19~4_combout  & (((!\Mux19~5_combout ))))

	.dataa(\Mux19~8_combout ),
	.datab(\ShiftRight0~108_combout ),
	.datac(\Mux19~4_combout ),
	.datad(\Mux19~5_combout ),
	.cin(gnd),
	.combout(\Mux19~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~9 .lut_mask = 16'hC0AF;
defparam \Mux19~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y43_N4
cycloneive_lcell_comb \Mux19~10 (
// Equation(s):
// \Mux19~10_combout  = (\Mux19~3_combout  & (((\Mux19~9_combout )))) # (!\Mux19~3_combout  & ((\Mux19~9_combout  & (\ShiftRight0~93_combout )) # (!\Mux19~9_combout  & ((\ShiftRight0~94_combout )))))

	.dataa(\ShiftRight0~93_combout ),
	.datab(\ShiftRight0~94_combout ),
	.datac(\Mux19~3_combout ),
	.datad(\Mux19~9_combout ),
	.cin(gnd),
	.combout(\Mux19~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~10 .lut_mask = 16'hFA0C;
defparam \Mux19~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N8
cycloneive_lcell_comb \Mux16~4 (
// Equation(s):
// \Mux16~4_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!Mux161 & !alu_a_mux_output_15)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (Mux161 $ (alu_a_mux_output_15))))

	.dataa(Mux161),
	.datab(alu_a_mux_output_15),
	.datac(\Mux19~2_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~4 .lut_mask = 16'hF016;
defparam \Mux16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N14
cycloneive_lcell_comb \Add0~51 (
// Equation(s):
// \Add0~51_combout  = Mux161 $ (temp_ALUop_output_0)

	.dataa(Mux161),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_ALUop_output_0),
	.cin(gnd),
	.combout(\Add0~51_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~51 .lut_mask = 16'h55AA;
defparam \Add0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N14
cycloneive_lcell_comb \Add0~53 (
// Equation(s):
// \Add0~53_combout  = (\Add0~52_combout  & ((alu_a_mux_output_14 & (\Add0~50  & VCC)) # (!alu_a_mux_output_14 & (!\Add0~50 )))) # (!\Add0~52_combout  & ((alu_a_mux_output_14 & (!\Add0~50 )) # (!alu_a_mux_output_14 & ((\Add0~50 ) # (GND)))))
// \Add0~54  = CARRY((\Add0~52_combout  & (!alu_a_mux_output_14 & !\Add0~50 )) # (!\Add0~52_combout  & ((!\Add0~50 ) # (!alu_a_mux_output_14))))

	.dataa(\Add0~52_combout ),
	.datab(alu_a_mux_output_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~50 ),
	.combout(\Add0~53_combout ),
	.cout(\Add0~54 ));
// synopsys translate_off
defparam \Add0~53 .lut_mask = 16'h9617;
defparam \Add0~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N16
cycloneive_lcell_comb \Add0~55 (
// Equation(s):
// \Add0~55_combout  = ((alu_a_mux_output_15 $ (\Add0~51_combout  $ (!\Add0~54 )))) # (GND)
// \Add0~56  = CARRY((alu_a_mux_output_15 & ((\Add0~51_combout ) # (!\Add0~54 ))) # (!alu_a_mux_output_15 & (\Add0~51_combout  & !\Add0~54 )))

	.dataa(alu_a_mux_output_15),
	.datab(\Add0~51_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~54 ),
	.combout(\Add0~55_combout ),
	.cout(\Add0~56 ));
// synopsys translate_off
defparam \Add0~55 .lut_mask = 16'h698E;
defparam \Add0~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N30
cycloneive_lcell_comb \ShiftLeft0~47 (
// Equation(s):
// \ShiftLeft0~47_combout  = (Mux301 & (alu_a_mux_output_9)) # (!Mux301 & ((alu_a_mux_output_11)))

	.dataa(gnd),
	.datab(alu_a_mux_output_9),
	.datac(alu_a_mux_output_11),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftLeft0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~47 .lut_mask = 16'hCCF0;
defparam \ShiftLeft0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N20
cycloneive_lcell_comb \ShiftLeft0~48 (
// Equation(s):
// \ShiftLeft0~48_combout  = (Mux311 & ((\ShiftLeft0~46_combout ))) # (!Mux311 & (\ShiftLeft0~47_combout ))

	.dataa(gnd),
	.datab(Mux311),
	.datac(\ShiftLeft0~47_combout ),
	.datad(\ShiftLeft0~46_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~48 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N22
cycloneive_lcell_comb \ShiftLeft0~65 (
// Equation(s):
// \ShiftLeft0~65_combout  = (Mux291 & ((\ShiftLeft0~48_combout ))) # (!Mux291 & (\ShiftLeft0~64_combout ))

	.dataa(\ShiftLeft0~64_combout ),
	.datab(gnd),
	.datac(Mux291),
	.datad(\ShiftLeft0~48_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~65 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N18
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (\Mux19~0_combout  & ((Mux281 & (\ShiftLeft0~34_combout )) # (!Mux281 & ((\ShiftLeft0~65_combout )))))

	.dataa(\ShiftLeft0~34_combout ),
	.datab(Mux281),
	.datac(\Mux19~0_combout ),
	.datad(\ShiftLeft0~65_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hB080;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N22
cycloneive_lcell_comb \Mux16~2 (
// Equation(s):
// \Mux16~2_combout  = (\Mux19~5_combout  & (\ShiftRight0~109_combout  & ((\Mux19~4_combout )))) # (!\Mux19~5_combout  & (((\Mux16~1_combout ) # (!\Mux19~4_combout ))))

	.dataa(\ShiftRight0~109_combout ),
	.datab(\Mux16~1_combout ),
	.datac(\Mux19~5_combout ),
	.datad(\Mux19~4_combout ),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~2 .lut_mask = 16'hAC0F;
defparam \Mux16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N10
cycloneive_lcell_comb \ShiftRight0~96 (
// Equation(s):
// \ShiftRight0~96_combout  = (Mux291 & (\ShiftRight0~87_combout )) # (!Mux291 & (((\ShiftRight0~77_combout ) # (\ShiftRight0~78_combout ))))

	.dataa(Mux291),
	.datab(\ShiftRight0~87_combout ),
	.datac(\ShiftRight0~77_combout ),
	.datad(\ShiftRight0~78_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~96 .lut_mask = 16'hDDD8;
defparam \ShiftRight0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N4
cycloneive_lcell_comb \Mux16~3 (
// Equation(s):
// \Mux16~3_combout  = (\Mux19~3_combout  & (((\Mux16~2_combout )))) # (!\Mux19~3_combout  & ((\Mux16~2_combout  & ((\ShiftRight0~96_combout ))) # (!\Mux16~2_combout  & (\ShiftRight0~97_combout ))))

	.dataa(\ShiftRight0~97_combout ),
	.datab(\Mux19~3_combout ),
	.datac(\Mux16~2_combout ),
	.datad(\ShiftRight0~96_combout ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~3 .lut_mask = 16'hF2C2;
defparam \Mux16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N2
cycloneive_lcell_comb \Add0~52 (
// Equation(s):
// \Add0~52_combout  = temp_ALUop_output_0 $ (((Mux17) # ((alu_b_mux_output_14 & !Mux16))))

	.dataa(temp_ALUop_output_0),
	.datab(alu_b_mux_output_14),
	.datac(Mux16),
	.datad(Mux17),
	.cin(gnd),
	.combout(\Add0~52_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~52 .lut_mask = 16'h55A6;
defparam \Add0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N8
cycloneive_lcell_comb \Mux17~4 (
// Equation(s):
// \Mux17~4_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!Mux171 & !alu_a_mux_output_14)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (Mux171 $ (alu_a_mux_output_14))))

	.dataa(Mux171),
	.datab(\Mux19~2_combout ),
	.datac(\Mux19~1_combout ),
	.datad(alu_a_mux_output_14),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~4 .lut_mask = 16'hC1C6;
defparam \Mux17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N18
cycloneive_lcell_comb \ShiftRight0~110 (
// Equation(s):
// \ShiftRight0~110_combout  = (!\ShiftLeft0~13_combout  & (!Mux281 & \ShiftRight0~44_combout ))

	.dataa(\ShiftLeft0~13_combout ),
	.datab(Mux281),
	.datac(\ShiftRight0~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~110_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~110 .lut_mask = 16'h1010;
defparam \ShiftRight0~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N18
cycloneive_lcell_comb \ShiftLeft0~62 (
// Equation(s):
// \ShiftLeft0~62_combout  = (Mux301 & ((alu_a_mux_output_12))) # (!Mux301 & (alu_a_mux_output_14))

	.dataa(Mux301),
	.datab(alu_a_mux_output_14),
	.datac(gnd),
	.datad(alu_a_mux_output_12),
	.cin(gnd),
	.combout(\ShiftLeft0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~62 .lut_mask = 16'hEE44;
defparam \ShiftLeft0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N12
cycloneive_lcell_comb \ShiftLeft0~66 (
// Equation(s):
// \ShiftLeft0~66_combout  = (Mux311 & (\ShiftLeft0~55_combout )) # (!Mux311 & ((\ShiftLeft0~62_combout )))

	.dataa(gnd),
	.datab(Mux311),
	.datac(\ShiftLeft0~55_combout ),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~66 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N12
cycloneive_lcell_comb \ShiftLeft0~67 (
// Equation(s):
// \ShiftLeft0~67_combout  = (Mux291 & (\ShiftLeft0~51_combout )) # (!Mux291 & ((\ShiftLeft0~66_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~51_combout ),
	.datac(Mux291),
	.datad(\ShiftLeft0~66_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~67 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N8
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (\Mux19~0_combout  & ((Mux281 & ((\ShiftLeft0~36_combout ))) # (!Mux281 & (\ShiftLeft0~67_combout ))))

	.dataa(\Mux19~0_combout ),
	.datab(\ShiftLeft0~67_combout ),
	.datac(Mux281),
	.datad(\ShiftLeft0~36_combout ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hA808;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N12
cycloneive_lcell_comb \Mux17~2 (
// Equation(s):
// \Mux17~2_combout  = (\Mux19~5_combout  & (\ShiftRight0~110_combout  & (\Mux19~4_combout ))) # (!\Mux19~5_combout  & (((\Mux17~1_combout ) # (!\Mux19~4_combout ))))

	.dataa(\Mux19~5_combout ),
	.datab(\ShiftRight0~110_combout ),
	.datac(\Mux19~4_combout ),
	.datad(\Mux17~1_combout ),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~2 .lut_mask = 16'hD585;
defparam \Mux17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N2
cycloneive_lcell_comb \Mux17~3 (
// Equation(s):
// \Mux17~3_combout  = (\Mux17~2_combout  & ((\Mux19~3_combout ) # ((\ShiftRight0~100_combout )))) # (!\Mux17~2_combout  & (!\Mux19~3_combout  & ((\ShiftRight0~101_combout ))))

	.dataa(\Mux17~2_combout ),
	.datab(\Mux19~3_combout ),
	.datac(\ShiftRight0~100_combout ),
	.datad(\ShiftRight0~101_combout ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~3 .lut_mask = 16'hB9A8;
defparam \Mux17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N18
cycloneive_lcell_comb \ShiftLeft0~70 (
// Equation(s):
// \ShiftLeft0~70_combout  = (Mux291 & ((\ShiftLeft0~56_combout ))) # (!Mux291 & (\ShiftLeft0~69_combout ))

	.dataa(\ShiftLeft0~69_combout ),
	.datab(gnd),
	.datac(Mux291),
	.datad(\ShiftLeft0~56_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~70 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N2
cycloneive_lcell_comb \Mux12~2 (
// Equation(s):
// \Mux12~2_combout  = (temp_ALUop_output_0) # ((\Mux19~0_combout  & Mux281))

	.dataa(temp_ALUop_output_0),
	.datab(gnd),
	.datac(\Mux19~0_combout ),
	.datad(Mux281),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~2 .lut_mask = 16'hFAAA;
defparam \Mux12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N24
cycloneive_lcell_comb \ShiftRight0~21 (
// Equation(s):
// \ShiftRight0~21_combout  = (Mux281 & ((Mux291 & (\ShiftRight0~18_combout )) # (!Mux291 & ((\ShiftRight0~20_combout )))))

	.dataa(\ShiftRight0~18_combout ),
	.datab(Mux291),
	.datac(\ShiftRight0~20_combout ),
	.datad(Mux281),
	.cin(gnd),
	.combout(\ShiftRight0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~21 .lut_mask = 16'hB800;
defparam \ShiftRight0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N28
cycloneive_lcell_comb \ShiftRight0~28 (
// Equation(s):
// \ShiftRight0~28_combout  = (\ShiftRight0~21_combout ) # ((!Mux281 & \ShiftRight0~27_combout ))

	.dataa(gnd),
	.datab(Mux281),
	.datac(\ShiftRight0~27_combout ),
	.datad(\ShiftRight0~21_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~28 .lut_mask = 16'hFF30;
defparam \ShiftRight0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N28
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (\Mux12~1_combout  & ((\Mux12~2_combout  & ((\ShiftRight0~28_combout ))) # (!\Mux12~2_combout  & (\ShiftLeft0~14_combout )))) # (!\Mux12~1_combout  & (((!\Mux12~2_combout ))))

	.dataa(\Mux12~1_combout ),
	.datab(\ShiftLeft0~14_combout ),
	.datac(\Mux12~2_combout ),
	.datad(\ShiftRight0~28_combout ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hAD0D;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N8
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (temp_ALUop_output_0) # ((\ShiftLeft0~10_combout ) # ((\ShiftLeft0~26_combout ) # (Mux271)))

	.dataa(temp_ALUop_output_0),
	.datab(\ShiftLeft0~10_combout ),
	.datac(\ShiftLeft0~26_combout ),
	.datad(Mux271),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hFFFE;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N16
cycloneive_lcell_comb \Mux14~2 (
// Equation(s):
// \Mux14~2_combout  = (\Mux14~1_combout  & ((\ShiftLeft0~70_combout ) # ((\Mux12~0_combout )))) # (!\Mux14~1_combout  & (((\ShiftLeft0~40_combout  & !\Mux12~0_combout ))))

	.dataa(\ShiftLeft0~70_combout ),
	.datab(\ShiftLeft0~40_combout ),
	.datac(\Mux14~1_combout ),
	.datad(\Mux12~0_combout ),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~2 .lut_mask = 16'hF0AC;
defparam \Mux14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N22
cycloneive_lcell_comb \Mux14~3 (
// Equation(s):
// \Mux14~3_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!alu_a_mux_output_17 & !Mux14)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (alu_a_mux_output_17 $ (Mux14))))

	.dataa(\Mux19~2_combout ),
	.datab(alu_a_mux_output_17),
	.datac(Mux14),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~3 .lut_mask = 16'hAA16;
defparam \Mux14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N8
cycloneive_lcell_comb \Add0~57 (
// Equation(s):
// \Add0~57_combout  = Mux14 $ (temp_ALUop_output_0)

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux14),
	.datad(temp_ALUop_output_0),
	.cin(gnd),
	.combout(\Add0~57_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~57 .lut_mask = 16'h0FF0;
defparam \Add0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N18
cycloneive_lcell_comb \Add0~59 (
// Equation(s):
// \Add0~59_combout  = (\Add0~58_combout  & ((alu_a_mux_output_16 & (\Add0~56  & VCC)) # (!alu_a_mux_output_16 & (!\Add0~56 )))) # (!\Add0~58_combout  & ((alu_a_mux_output_16 & (!\Add0~56 )) # (!alu_a_mux_output_16 & ((\Add0~56 ) # (GND)))))
// \Add0~60  = CARRY((\Add0~58_combout  & (!alu_a_mux_output_16 & !\Add0~56 )) # (!\Add0~58_combout  & ((!\Add0~56 ) # (!alu_a_mux_output_16))))

	.dataa(\Add0~58_combout ),
	.datab(alu_a_mux_output_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~56 ),
	.combout(\Add0~59_combout ),
	.cout(\Add0~60 ));
// synopsys translate_off
defparam \Add0~59 .lut_mask = 16'h9617;
defparam \Add0~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N20
cycloneive_lcell_comb \Add0~61 (
// Equation(s):
// \Add0~61_combout  = ((alu_a_mux_output_17 $ (\Add0~57_combout  $ (!\Add0~60 )))) # (GND)
// \Add0~62  = CARRY((alu_a_mux_output_17 & ((\Add0~57_combout ) # (!\Add0~60 ))) # (!alu_a_mux_output_17 & (\Add0~57_combout  & !\Add0~60 )))

	.dataa(alu_a_mux_output_17),
	.datab(\Add0~57_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~60 ),
	.combout(\Add0~61_combout ),
	.cout(\Add0~62 ));
// synopsys translate_off
defparam \Add0~61 .lut_mask = 16'h698E;
defparam \Add0~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N6
cycloneive_lcell_comb \Add0~58 (
// Equation(s):
// \Add0~58_combout  = Mux15 $ (temp_ALUop_output_0)

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux15),
	.datad(temp_ALUop_output_0),
	.cin(gnd),
	.combout(\Add0~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~58 .lut_mask = 16'h0FF0;
defparam \Add0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N4
cycloneive_lcell_comb \ShiftRight0~55 (
// Equation(s):
// \ShiftRight0~55_combout  = (\ShiftRight0~52_combout ) # ((Mux281 & (!Mux291 & \ShiftRight0~54_combout )))

	.dataa(\ShiftRight0~52_combout ),
	.datab(Mux281),
	.datac(Mux291),
	.datad(\ShiftRight0~54_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~55 .lut_mask = 16'hAEAA;
defparam \ShiftRight0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N20
cycloneive_lcell_comb \ShiftLeft0~17 (
// Equation(s):
// \ShiftLeft0~17_combout  = (\ShiftLeft0~16_combout  & (!Mux291 & (!\ShiftLeft0~11_combout  & !Mux281)))

	.dataa(\ShiftLeft0~16_combout ),
	.datab(Mux291),
	.datac(\ShiftLeft0~11_combout ),
	.datad(Mux281),
	.cin(gnd),
	.combout(\ShiftLeft0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~17 .lut_mask = 16'h0002;
defparam \ShiftLeft0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N2
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (\Mux12~1_combout  & ((\Mux12~2_combout  & (\ShiftRight0~55_combout )) # (!\Mux12~2_combout  & ((\ShiftLeft0~17_combout ))))) # (!\Mux12~1_combout  & (((!\Mux12~2_combout ))))

	.dataa(\Mux12~1_combout ),
	.datab(\ShiftRight0~55_combout ),
	.datac(\Mux12~2_combout ),
	.datad(\ShiftLeft0~17_combout ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'h8F85;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N24
cycloneive_lcell_comb \ShiftLeft0~59 (
// Equation(s):
// \ShiftLeft0~59_combout  = (Mux311 & (\ShiftLeft0~47_combout )) # (!Mux311 & ((\ShiftLeft0~54_combout )))

	.dataa(gnd),
	.datab(Mux311),
	.datac(\ShiftLeft0~47_combout ),
	.datad(\ShiftLeft0~54_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~59 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y41_N18
cycloneive_lcell_comb \ShiftLeft0~72 (
// Equation(s):
// \ShiftLeft0~72_combout  = (!Mux311 & ((Mux301 & (alu_a_mux_output_14)) # (!Mux301 & ((alu_a_mux_output_16)))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_14),
	.datac(Mux311),
	.datad(alu_a_mux_output_16),
	.cin(gnd),
	.combout(\ShiftLeft0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~72 .lut_mask = 16'h0D08;
defparam \ShiftLeft0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N30
cycloneive_lcell_comb \ShiftLeft0~73 (
// Equation(s):
// \ShiftLeft0~73_combout  = (Mux291 & (((\ShiftLeft0~59_combout )))) # (!Mux291 & ((\ShiftLeft0~71_combout ) # ((\ShiftLeft0~72_combout ))))

	.dataa(\ShiftLeft0~71_combout ),
	.datab(\ShiftLeft0~59_combout ),
	.datac(Mux291),
	.datad(\ShiftLeft0~72_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~73 .lut_mask = 16'hCFCA;
defparam \ShiftLeft0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N16
cycloneive_lcell_comb \Mux15~2 (
// Equation(s):
// \Mux15~2_combout  = (\Mux15~1_combout  & (((\ShiftLeft0~73_combout ) # (\Mux12~0_combout )))) # (!\Mux15~1_combout  & (\ShiftLeft0~44_combout  & ((!\Mux12~0_combout ))))

	.dataa(\ShiftLeft0~44_combout ),
	.datab(\Mux15~1_combout ),
	.datac(\ShiftLeft0~73_combout ),
	.datad(\Mux12~0_combout ),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~2 .lut_mask = 16'hCCE2;
defparam \Mux15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N2
cycloneive_lcell_comb \Mux15~3 (
// Equation(s):
// \Mux15~3_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!Mux15 & !alu_a_mux_output_16)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (Mux15 $ (alu_a_mux_output_16))))

	.dataa(\Mux19~2_combout ),
	.datab(Mux15),
	.datac(\Mux19~1_combout ),
	.datad(alu_a_mux_output_16),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~3 .lut_mask = 16'hA1A6;
defparam \Mux15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N30
cycloneive_lcell_comb \Add0~63 (
// Equation(s):
// \Add0~63_combout  = temp_ALUop_output_0 $ (Mux12)

	.dataa(gnd),
	.datab(temp_ALUop_output_0),
	.datac(gnd),
	.datad(Mux12),
	.cin(gnd),
	.combout(\Add0~63_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~63 .lut_mask = 16'h33CC;
defparam \Add0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N22
cycloneive_lcell_comb \Add0~65 (
// Equation(s):
// \Add0~65_combout  = (\Add0~64_combout  & ((alu_a_mux_output_18 & (\Add0~62  & VCC)) # (!alu_a_mux_output_18 & (!\Add0~62 )))) # (!\Add0~64_combout  & ((alu_a_mux_output_18 & (!\Add0~62 )) # (!alu_a_mux_output_18 & ((\Add0~62 ) # (GND)))))
// \Add0~66  = CARRY((\Add0~64_combout  & (!alu_a_mux_output_18 & !\Add0~62 )) # (!\Add0~64_combout  & ((!\Add0~62 ) # (!alu_a_mux_output_18))))

	.dataa(\Add0~64_combout ),
	.datab(alu_a_mux_output_18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~62 ),
	.combout(\Add0~65_combout ),
	.cout(\Add0~66 ));
// synopsys translate_off
defparam \Add0~65 .lut_mask = 16'h9617;
defparam \Add0~65 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N24
cycloneive_lcell_comb \Add0~67 (
// Equation(s):
// \Add0~67_combout  = ((\Add0~63_combout  $ (alu_a_mux_output_19 $ (!\Add0~66 )))) # (GND)
// \Add0~68  = CARRY((\Add0~63_combout  & ((alu_a_mux_output_19) # (!\Add0~66 ))) # (!\Add0~63_combout  & (alu_a_mux_output_19 & !\Add0~66 )))

	.dataa(\Add0~63_combout ),
	.datab(alu_a_mux_output_19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~66 ),
	.combout(\Add0~67_combout ),
	.cout(\Add0~68 ));
// synopsys translate_off
defparam \Add0~67 .lut_mask = 16'h698E;
defparam \Add0~67 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N30
cycloneive_lcell_comb \ShiftLeft0~49 (
// Equation(s):
// \ShiftLeft0~49_combout  = (Mux291 & (\ShiftLeft0~33_combout )) # (!Mux291 & ((\ShiftLeft0~48_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~33_combout ),
	.datac(Mux291),
	.datad(\ShiftLeft0~48_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~49 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N30
cycloneive_lcell_comb \ShiftLeft0~74 (
// Equation(s):
// \ShiftLeft0~74_combout  = (Mux311 & ((Mux301 & ((alu_a_mux_output_16))) # (!Mux301 & (alu_a_mux_output_18))))

	.dataa(alu_a_mux_output_18),
	.datab(Mux311),
	.datac(Mux301),
	.datad(alu_a_mux_output_16),
	.cin(gnd),
	.combout(\ShiftLeft0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~74 .lut_mask = 16'hC808;
defparam \ShiftLeft0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N4
cycloneive_lcell_comb \ShiftLeft0~63 (
// Equation(s):
// \ShiftLeft0~63_combout  = (Mux301 & ((alu_a_mux_output_13))) # (!Mux301 & (alu_a_mux_output_15))

	.dataa(alu_a_mux_output_15),
	.datab(gnd),
	.datac(alu_a_mux_output_13),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftLeft0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~63 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N26
cycloneive_lcell_comb \ShiftLeft0~64 (
// Equation(s):
// \ShiftLeft0~64_combout  = (Mux311 & ((\ShiftLeft0~62_combout ))) # (!Mux311 & (\ShiftLeft0~63_combout ))

	.dataa(gnd),
	.datab(Mux311),
	.datac(\ShiftLeft0~63_combout ),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~64 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N28
cycloneive_lcell_comb \ShiftLeft0~76 (
// Equation(s):
// \ShiftLeft0~76_combout  = (Mux291 & (((\ShiftLeft0~64_combout )))) # (!Mux291 & ((\ShiftLeft0~75_combout ) # ((\ShiftLeft0~74_combout ))))

	.dataa(\ShiftLeft0~75_combout ),
	.datab(Mux291),
	.datac(\ShiftLeft0~74_combout ),
	.datad(\ShiftLeft0~64_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~76 .lut_mask = 16'hFE32;
defparam \ShiftLeft0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N24
cycloneive_lcell_comb \ShiftRight0~89 (
// Equation(s):
// \ShiftRight0~89_combout  = (Mux281 & ((\ShiftRight0~83_combout ))) # (!Mux281 & (\ShiftRight0~88_combout ))

	.dataa(\ShiftRight0~88_combout ),
	.datab(gnd),
	.datac(Mux281),
	.datad(\ShiftRight0~83_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~89 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N30
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = temp_ALUop_output_0 $ (!\Mux19~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(\Mux19~0_combout ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hF00F;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N24
cycloneive_lcell_comb \Mux12~5 (
// Equation(s):
// \Mux12~5_combout  = (\Mux12~2_combout  & (((\ShiftRight0~89_combout  & \Mux12~1_combout )))) # (!\Mux12~2_combout  & ((\Mux12~4_combout ) # ((!\Mux12~1_combout ))))

	.dataa(\Mux12~4_combout ),
	.datab(\ShiftRight0~89_combout ),
	.datac(\Mux12~2_combout ),
	.datad(\Mux12~1_combout ),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~5 .lut_mask = 16'hCA0F;
defparam \Mux12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N6
cycloneive_lcell_comb \Mux12~6 (
// Equation(s):
// \Mux12~6_combout  = (\Mux12~0_combout  & (((\Mux12~5_combout )))) # (!\Mux12~0_combout  & ((\Mux12~5_combout  & ((\ShiftLeft0~76_combout ))) # (!\Mux12~5_combout  & (\ShiftLeft0~49_combout ))))

	.dataa(\ShiftLeft0~49_combout ),
	.datab(\ShiftLeft0~76_combout ),
	.datac(\Mux12~0_combout ),
	.datad(\Mux12~5_combout ),
	.cin(gnd),
	.combout(\Mux12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~6 .lut_mask = 16'hFC0A;
defparam \Mux12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y42_N24
cycloneive_lcell_comb \Mux12~7 (
// Equation(s):
// \Mux12~7_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!alu_a_mux_output_19 & !Mux12)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (alu_a_mux_output_19 $ (Mux12))))

	.dataa(alu_a_mux_output_19),
	.datab(Mux12),
	.datac(\Mux19~2_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~7 .lut_mask = 16'hF016;
defparam \Mux12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N28
cycloneive_lcell_comb \Mux13~4 (
// Equation(s):
// \Mux13~4_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!alu_a_mux_output_18 & !Mux13)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (alu_a_mux_output_18 $ (Mux13))))

	.dataa(\Mux19~2_combout ),
	.datab(alu_a_mux_output_18),
	.datac(Mux13),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~4 .lut_mask = 16'hAA16;
defparam \Mux13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N24
cycloneive_lcell_comb \ShiftLeft0~78 (
// Equation(s):
// \ShiftLeft0~78_combout  = (!Mux311 & ((Mux301 & ((alu_a_mux_output_16))) # (!Mux301 & (alu_a_mux_output_18))))

	.dataa(alu_a_mux_output_18),
	.datab(Mux311),
	.datac(Mux301),
	.datad(alu_a_mux_output_16),
	.cin(gnd),
	.combout(\ShiftLeft0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~78 .lut_mask = 16'h3202;
defparam \ShiftLeft0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N14
cycloneive_lcell_comb \ShiftLeft0~77 (
// Equation(s):
// \ShiftLeft0~77_combout  = (Mux311 & ((Mux301 & ((alu_a_mux_output_15))) # (!Mux301 & (alu_a_mux_output_17))))

	.dataa(alu_a_mux_output_17),
	.datab(Mux301),
	.datac(Mux311),
	.datad(alu_a_mux_output_15),
	.cin(gnd),
	.combout(\ShiftLeft0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~77 .lut_mask = 16'hE020;
defparam \ShiftLeft0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N24
cycloneive_lcell_comb \ShiftLeft0~79 (
// Equation(s):
// \ShiftLeft0~79_combout  = (Mux291 & (((\ShiftLeft0~66_combout )))) # (!Mux291 & ((\ShiftLeft0~78_combout ) # ((\ShiftLeft0~77_combout ))))

	.dataa(Mux291),
	.datab(\ShiftLeft0~78_combout ),
	.datac(\ShiftLeft0~77_combout ),
	.datad(\ShiftLeft0~66_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~79 .lut_mask = 16'hFE54;
defparam \ShiftLeft0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N22
cycloneive_lcell_comb \Mux13~2 (
// Equation(s):
// \Mux13~2_combout  = (\Mux12~1_combout  & ((\Mux12~2_combout  & ((\ShiftRight0~74_combout ))) # (!\Mux12~2_combout  & (\Mux13~1_combout )))) # (!\Mux12~1_combout  & (((!\Mux12~2_combout ))))

	.dataa(\Mux13~1_combout ),
	.datab(\Mux12~1_combout ),
	.datac(\Mux12~2_combout ),
	.datad(\ShiftRight0~74_combout ),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~2 .lut_mask = 16'hCB0B;
defparam \Mux13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N26
cycloneive_lcell_comb \Mux13~3 (
// Equation(s):
// \Mux13~3_combout  = (\Mux12~0_combout  & (((\Mux13~2_combout )))) # (!\Mux12~0_combout  & ((\Mux13~2_combout  & ((\ShiftLeft0~79_combout ))) # (!\Mux13~2_combout  & (\ShiftLeft0~52_combout ))))

	.dataa(\ShiftLeft0~52_combout ),
	.datab(\Mux12~0_combout ),
	.datac(\ShiftLeft0~79_combout ),
	.datad(\Mux13~2_combout ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~3 .lut_mask = 16'hFC22;
defparam \Mux13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N4
cycloneive_lcell_comb \Add0~64 (
// Equation(s):
// \Add0~64_combout  = Mux13 $ (temp_ALUop_output_0)

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux13),
	.datad(temp_ALUop_output_0),
	.cin(gnd),
	.combout(\Add0~64_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~64 .lut_mask = 16'h0FF0;
defparam \Add0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N10
cycloneive_lcell_comb \ShiftLeft0~60 (
// Equation(s):
// \ShiftLeft0~60_combout  = (Mux291 & ((\ShiftLeft0~42_combout ) # ((\ShiftLeft0~43_combout )))) # (!Mux291 & (((\ShiftLeft0~59_combout ))))

	.dataa(\ShiftLeft0~42_combout ),
	.datab(\ShiftLeft0~59_combout ),
	.datac(Mux291),
	.datad(\ShiftLeft0~43_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~60 .lut_mask = 16'hFCAC;
defparam \ShiftLeft0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N24
cycloneive_lcell_comb \ShiftLeft0~80 (
// Equation(s):
// \ShiftLeft0~80_combout  = (Mux311 & (((Mux301)))) # (!Mux311 & ((Mux301 & (alu_a_mux_output_18)) # (!Mux301 & ((alu_a_mux_output_20)))))

	.dataa(Mux311),
	.datab(alu_a_mux_output_18),
	.datac(Mux301),
	.datad(alu_a_mux_output_20),
	.cin(gnd),
	.combout(\ShiftLeft0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~80 .lut_mask = 16'hE5E0;
defparam \ShiftLeft0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N30
cycloneive_lcell_comb \ShiftLeft0~81 (
// Equation(s):
// \ShiftLeft0~81_combout  = (Mux311 & ((\ShiftLeft0~80_combout  & (alu_a_mux_output_17)) # (!\ShiftLeft0~80_combout  & ((alu_a_mux_output_19))))) # (!Mux311 & (((\ShiftLeft0~80_combout ))))

	.dataa(alu_a_mux_output_17),
	.datab(alu_a_mux_output_19),
	.datac(Mux311),
	.datad(\ShiftLeft0~80_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~81 .lut_mask = 16'hAFC0;
defparam \ShiftLeft0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y39_N6
cycloneive_lcell_comb \ShiftLeft0~71 (
// Equation(s):
// \ShiftLeft0~71_combout  = (Mux311 & ((Mux301 & (alu_a_mux_output_13)) # (!Mux301 & ((alu_a_mux_output_15)))))

	.dataa(Mux301),
	.datab(Mux311),
	.datac(alu_a_mux_output_13),
	.datad(alu_a_mux_output_15),
	.cin(gnd),
	.combout(\ShiftLeft0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~71 .lut_mask = 16'hC480;
defparam \ShiftLeft0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N18
cycloneive_lcell_comb \ShiftLeft0~82 (
// Equation(s):
// \ShiftLeft0~82_combout  = (Mux291 & ((\ShiftLeft0~72_combout ) # ((\ShiftLeft0~71_combout )))) # (!Mux291 & (((\ShiftLeft0~81_combout ))))

	.dataa(Mux291),
	.datab(\ShiftLeft0~72_combout ),
	.datac(\ShiftLeft0~81_combout ),
	.datad(\ShiftLeft0~71_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~82 .lut_mask = 16'hFAD8;
defparam \ShiftLeft0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y41_N14
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (!Mux281 & (!\ShiftLeft0~26_combout  & (\ShiftLeft0~29_combout  & !\ShiftLeft0~10_combout )))

	.dataa(Mux281),
	.datab(\ShiftLeft0~26_combout ),
	.datac(\ShiftLeft0~29_combout ),
	.datad(\ShiftLeft0~10_combout ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'h0010;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N16
cycloneive_lcell_comb \Mux11~2 (
// Equation(s):
// \Mux11~2_combout  = (\Mux12~1_combout  & ((\Mux12~2_combout  & ((\ShiftRight0~95_combout ))) # (!\Mux12~2_combout  & (\Mux11~1_combout )))) # (!\Mux12~1_combout  & (((!\Mux12~2_combout ))))

	.dataa(\Mux12~1_combout ),
	.datab(\Mux11~1_combout ),
	.datac(\Mux12~2_combout ),
	.datad(\ShiftRight0~95_combout ),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~2 .lut_mask = 16'hAD0D;
defparam \Mux11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N28
cycloneive_lcell_comb \Mux11~3 (
// Equation(s):
// \Mux11~3_combout  = (\Mux12~0_combout  & (((\Mux11~2_combout )))) # (!\Mux12~0_combout  & ((\Mux11~2_combout  & ((\ShiftLeft0~82_combout ))) # (!\Mux11~2_combout  & (\ShiftLeft0~60_combout ))))

	.dataa(\ShiftLeft0~60_combout ),
	.datab(\ShiftLeft0~82_combout ),
	.datac(\Mux12~0_combout ),
	.datad(\Mux11~2_combout ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~3 .lut_mask = 16'hFC0A;
defparam \Mux11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N0
cycloneive_lcell_comb \Add0~69 (
// Equation(s):
// \Add0~69_combout  = Mux11 $ (temp_ALUop_output_0)

	.dataa(gnd),
	.datab(Mux11),
	.datac(temp_ALUop_output_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add0~69_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~69 .lut_mask = 16'h3C3C;
defparam \Add0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N26
cycloneive_lcell_comb \Add0~70 (
// Equation(s):
// \Add0~70_combout  = (alu_a_mux_output_20 & ((\Add0~69_combout  & (\Add0~68  & VCC)) # (!\Add0~69_combout  & (!\Add0~68 )))) # (!alu_a_mux_output_20 & ((\Add0~69_combout  & (!\Add0~68 )) # (!\Add0~69_combout  & ((\Add0~68 ) # (GND)))))
// \Add0~71  = CARRY((alu_a_mux_output_20 & (!\Add0~69_combout  & !\Add0~68 )) # (!alu_a_mux_output_20 & ((!\Add0~68 ) # (!\Add0~69_combout ))))

	.dataa(alu_a_mux_output_20),
	.datab(\Add0~69_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~68 ),
	.combout(\Add0~70_combout ),
	.cout(\Add0~71 ));
// synopsys translate_off
defparam \Add0~70 .lut_mask = 16'h9617;
defparam \Add0~70 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X68_Y43_N2
cycloneive_lcell_comb \Mux11~4 (
// Equation(s):
// \Mux11~4_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!alu_a_mux_output_20 & !Mux11)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (alu_a_mux_output_20 $ (Mux11))))

	.dataa(alu_a_mux_output_20),
	.datab(\Mux19~2_combout ),
	.datac(\Mux19~1_combout ),
	.datad(Mux11),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~4 .lut_mask = 16'hC1C6;
defparam \Mux11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N26
cycloneive_lcell_comb \Add0~72 (
// Equation(s):
// \Add0~72_combout  = temp_ALUop_output_0 $ (Mux10)

	.dataa(gnd),
	.datab(temp_ALUop_output_0),
	.datac(gnd),
	.datad(Mux10),
	.cin(gnd),
	.combout(\Add0~72_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~72 .lut_mask = 16'h33CC;
defparam \Add0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N28
cycloneive_lcell_comb \Add0~73 (
// Equation(s):
// \Add0~73_combout  = ((alu_a_mux_output_21 $ (\Add0~72_combout  $ (!\Add0~71 )))) # (GND)
// \Add0~74  = CARRY((alu_a_mux_output_21 & ((\Add0~72_combout ) # (!\Add0~71 ))) # (!alu_a_mux_output_21 & (\Add0~72_combout  & !\Add0~71 )))

	.dataa(alu_a_mux_output_21),
	.datab(\Add0~72_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~71 ),
	.combout(\Add0~73_combout ),
	.cout(\Add0~74 ));
// synopsys translate_off
defparam \Add0~73 .lut_mask = 16'h698E;
defparam \Add0~73 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N26
cycloneive_lcell_comb \ShiftLeft0~83 (
// Equation(s):
// \ShiftLeft0~83_combout  = (Mux311 & (((Mux301)))) # (!Mux311 & ((Mux301 & ((alu_a_mux_output_19))) # (!Mux301 & (alu_a_mux_output_21))))

	.dataa(alu_a_mux_output_21),
	.datab(Mux311),
	.datac(Mux301),
	.datad(alu_a_mux_output_19),
	.cin(gnd),
	.combout(\ShiftLeft0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~83 .lut_mask = 16'hF2C2;
defparam \ShiftLeft0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N0
cycloneive_lcell_comb \ShiftLeft0~84 (
// Equation(s):
// \ShiftLeft0~84_combout  = (Mux311 & ((\ShiftLeft0~83_combout  & (alu_a_mux_output_18)) # (!\ShiftLeft0~83_combout  & ((alu_a_mux_output_20))))) # (!Mux311 & (((\ShiftLeft0~83_combout ))))

	.dataa(alu_a_mux_output_18),
	.datab(Mux311),
	.datac(\ShiftLeft0~83_combout ),
	.datad(alu_a_mux_output_20),
	.cin(gnd),
	.combout(\ShiftLeft0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~84 .lut_mask = 16'hBCB0;
defparam \ShiftLeft0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N22
cycloneive_lcell_comb \ShiftLeft0~68 (
// Equation(s):
// \ShiftLeft0~68_combout  = (Mux301 & ((Mux311 & (alu_a_mux_output_14)) # (!Mux311 & ((alu_a_mux_output_15)))))

	.dataa(Mux311),
	.datab(Mux301),
	.datac(alu_a_mux_output_14),
	.datad(alu_a_mux_output_15),
	.cin(gnd),
	.combout(\ShiftLeft0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~68 .lut_mask = 16'hC480;
defparam \ShiftLeft0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N6
cycloneive_lcell_comb \ShiftRight0~22 (
// Equation(s):
// \ShiftRight0~22_combout  = (!Mux311 & (!Mux301 & alu_a_mux_output_17))

	.dataa(Mux311),
	.datab(Mux301),
	.datac(gnd),
	.datad(alu_a_mux_output_17),
	.cin(gnd),
	.combout(\ShiftRight0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~22 .lut_mask = 16'h1100;
defparam \ShiftRight0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N20
cycloneive_lcell_comb \ShiftLeft0~69 (
// Equation(s):
// \ShiftLeft0~69_combout  = (\ShiftLeft0~68_combout ) # ((\ShiftRight0~22_combout ) # ((\Mux1~0_combout  & alu_a_mux_output_16)))

	.dataa(\Mux1~0_combout ),
	.datab(alu_a_mux_output_16),
	.datac(\ShiftLeft0~68_combout ),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~69 .lut_mask = 16'hFFF8;
defparam \ShiftLeft0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N18
cycloneive_lcell_comb \ShiftLeft0~85 (
// Equation(s):
// \ShiftLeft0~85_combout  = (Mux291 & ((\ShiftLeft0~69_combout ))) # (!Mux291 & (\ShiftLeft0~84_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~84_combout ),
	.datac(Mux291),
	.datad(\ShiftLeft0~69_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~85 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N12
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (!\ShiftLeft0~10_combout  & (!\ShiftLeft0~26_combout  & (!Mux281 & \ShiftLeft0~25_combout )))

	.dataa(\ShiftLeft0~10_combout ),
	.datab(\ShiftLeft0~26_combout ),
	.datac(Mux281),
	.datad(\ShiftLeft0~25_combout ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'h0100;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N30
cycloneive_lcell_comb \Mux10~2 (
// Equation(s):
// \Mux10~2_combout  = (\Mux12~2_combout  & (\ShiftRight0~92_combout  & (\Mux12~1_combout ))) # (!\Mux12~2_combout  & (((\Mux10~1_combout ) # (!\Mux12~1_combout ))))

	.dataa(\ShiftRight0~92_combout ),
	.datab(\Mux12~2_combout ),
	.datac(\Mux12~1_combout ),
	.datad(\Mux10~1_combout ),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~2 .lut_mask = 16'hB383;
defparam \Mux10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N4
cycloneive_lcell_comb \Mux10~3 (
// Equation(s):
// \Mux10~3_combout  = (\Mux12~0_combout  & (((\Mux10~2_combout )))) # (!\Mux12~0_combout  & ((\Mux10~2_combout  & ((\ShiftLeft0~85_combout ))) # (!\Mux10~2_combout  & (\ShiftLeft0~57_combout ))))

	.dataa(\ShiftLeft0~57_combout ),
	.datab(\ShiftLeft0~85_combout ),
	.datac(\Mux12~0_combout ),
	.datad(\Mux10~2_combout ),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~3 .lut_mask = 16'hFC0A;
defparam \Mux10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N24
cycloneive_lcell_comb \Mux10~4 (
// Equation(s):
// \Mux10~4_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!alu_a_mux_output_21 & !Mux10)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (alu_a_mux_output_21 $ (Mux10))))

	.dataa(alu_a_mux_output_21),
	.datab(Mux10),
	.datac(\Mux19~2_combout ),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~4 .lut_mask = 16'hF016;
defparam \Mux10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N14
cycloneive_lcell_comb \Mux8~4 (
// Equation(s):
// \Mux8~4_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!Mux8 & !alu_a_mux_output_23)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (Mux8 $ (alu_a_mux_output_23))))

	.dataa(\Mux19~2_combout ),
	.datab(\Mux19~1_combout ),
	.datac(Mux8),
	.datad(alu_a_mux_output_23),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~4 .lut_mask = 16'h899A;
defparam \Mux8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N16
cycloneive_lcell_comb \ShiftLeft0~86 (
// Equation(s):
// \ShiftLeft0~86_combout  = (Mux311 & (((Mux301)))) # (!Mux311 & ((Mux301 & (alu_a_mux_output_21)) # (!Mux301 & ((alu_a_mux_output_23)))))

	.dataa(Mux311),
	.datab(alu_a_mux_output_21),
	.datac(Mux301),
	.datad(alu_a_mux_output_23),
	.cin(gnd),
	.combout(\ShiftLeft0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~86 .lut_mask = 16'hE5E0;
defparam \ShiftLeft0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N30
cycloneive_lcell_comb \ShiftLeft0~87 (
// Equation(s):
// \ShiftLeft0~87_combout  = (Mux311 & ((\ShiftLeft0~86_combout  & ((alu_a_mux_output_20))) # (!\ShiftLeft0~86_combout  & (alu_a_mux_output_22)))) # (!Mux311 & (((\ShiftLeft0~86_combout ))))

	.dataa(Mux311),
	.datab(alu_a_mux_output_22),
	.datac(alu_a_mux_output_20),
	.datad(\ShiftLeft0~86_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~87 .lut_mask = 16'hF588;
defparam \ShiftLeft0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N26
cycloneive_lcell_comb \ShiftLeft0~88 (
// Equation(s):
// \ShiftLeft0~88_combout  = (Mux291 & ((\ShiftLeft0~75_combout ) # ((\ShiftLeft0~74_combout )))) # (!Mux291 & (((\ShiftLeft0~87_combout ))))

	.dataa(\ShiftLeft0~75_combout ),
	.datab(Mux291),
	.datac(\ShiftLeft0~74_combout ),
	.datad(\ShiftLeft0~87_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~88 .lut_mask = 16'hFBC8;
defparam \ShiftLeft0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N28
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (!\ShiftLeft0~10_combout  & (!\ShiftLeft0~26_combout  & (!Mux281 & \ShiftLeft0~34_combout )))

	.dataa(\ShiftLeft0~10_combout ),
	.datab(\ShiftLeft0~26_combout ),
	.datac(Mux281),
	.datad(\ShiftLeft0~34_combout ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'h0100;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N18
cycloneive_lcell_comb \Mux8~2 (
// Equation(s):
// \Mux8~2_combout  = (\Mux12~2_combout  & (\ShiftRight0~98_combout  & (\Mux12~1_combout ))) # (!\Mux12~2_combout  & (((\Mux8~1_combout ) # (!\Mux12~1_combout ))))

	.dataa(\ShiftRight0~98_combout ),
	.datab(\Mux12~2_combout ),
	.datac(\Mux12~1_combout ),
	.datad(\Mux8~1_combout ),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~2 .lut_mask = 16'hB383;
defparam \Mux8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y40_N22
cycloneive_lcell_comb \Mux8~3 (
// Equation(s):
// \Mux8~3_combout  = (\Mux12~0_combout  & (((\Mux8~2_combout )))) # (!\Mux12~0_combout  & ((\Mux8~2_combout  & (\ShiftLeft0~88_combout )) # (!\Mux8~2_combout  & ((\ShiftLeft0~65_combout )))))

	.dataa(\ShiftLeft0~88_combout ),
	.datab(\ShiftLeft0~65_combout ),
	.datac(\Mux12~0_combout ),
	.datad(\Mux8~2_combout ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~3 .lut_mask = 16'hFA0C;
defparam \Mux8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N20
cycloneive_lcell_comb \Add0~75 (
// Equation(s):
// \Add0~75_combout  = Mux8 $ (temp_ALUop_output_0)

	.dataa(gnd),
	.datab(Mux8),
	.datac(temp_ALUop_output_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add0~75_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~75 .lut_mask = 16'h3C3C;
defparam \Add0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N16
cycloneive_lcell_comb \Add0~76 (
// Equation(s):
// \Add0~76_combout  = temp_ALUop_output_0 $ (Mux9)

	.dataa(gnd),
	.datab(temp_ALUop_output_0),
	.datac(gnd),
	.datad(Mux9),
	.cin(gnd),
	.combout(\Add0~76_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~76 .lut_mask = 16'h33CC;
defparam \Add0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N30
cycloneive_lcell_comb \Add0~77 (
// Equation(s):
// \Add0~77_combout  = (alu_a_mux_output_22 & ((\Add0~76_combout  & (\Add0~74  & VCC)) # (!\Add0~76_combout  & (!\Add0~74 )))) # (!alu_a_mux_output_22 & ((\Add0~76_combout  & (!\Add0~74 )) # (!\Add0~76_combout  & ((\Add0~74 ) # (GND)))))
// \Add0~78  = CARRY((alu_a_mux_output_22 & (!\Add0~76_combout  & !\Add0~74 )) # (!alu_a_mux_output_22 & ((!\Add0~74 ) # (!\Add0~76_combout ))))

	.dataa(alu_a_mux_output_22),
	.datab(\Add0~76_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~74 ),
	.combout(\Add0~77_combout ),
	.cout(\Add0~78 ));
// synopsys translate_off
defparam \Add0~77 .lut_mask = 16'h9617;
defparam \Add0~77 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N0
cycloneive_lcell_comb \Add0~79 (
// Equation(s):
// \Add0~79_combout  = ((alu_a_mux_output_23 $ (\Add0~75_combout  $ (!\Add0~78 )))) # (GND)
// \Add0~80  = CARRY((alu_a_mux_output_23 & ((\Add0~75_combout ) # (!\Add0~78 ))) # (!alu_a_mux_output_23 & (\Add0~75_combout  & !\Add0~78 )))

	.dataa(alu_a_mux_output_23),
	.datab(\Add0~75_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~78 ),
	.combout(\Add0~79_combout ),
	.cout(\Add0~80 ));
// synopsys translate_off
defparam \Add0~79 .lut_mask = 16'h698E;
defparam \Add0~79 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N12
cycloneive_lcell_comb \Mux9~4 (
// Equation(s):
// \Mux9~4_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!Mux9 & !alu_a_mux_output_22)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (Mux9 $ (alu_a_mux_output_22))))

	.dataa(\Mux19~2_combout ),
	.datab(Mux9),
	.datac(alu_a_mux_output_22),
	.datad(\Mux19~1_combout ),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~4 .lut_mask = 16'hAA16;
defparam \Mux9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N28
cycloneive_lcell_comb \ShiftLeft0~89 (
// Equation(s):
// \ShiftLeft0~89_combout  = (Mux311 & ((Mux301 & (alu_a_mux_output_19)) # (!Mux301 & ((alu_a_mux_output_21))))) # (!Mux311 & (((Mux301))))

	.dataa(alu_a_mux_output_19),
	.datab(Mux311),
	.datac(Mux301),
	.datad(alu_a_mux_output_21),
	.cin(gnd),
	.combout(\ShiftLeft0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~89 .lut_mask = 16'hBCB0;
defparam \ShiftLeft0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N10
cycloneive_lcell_comb \ShiftLeft0~90 (
// Equation(s):
// \ShiftLeft0~90_combout  = (Mux311 & (((\ShiftLeft0~89_combout )))) # (!Mux311 & ((\ShiftLeft0~89_combout  & (alu_a_mux_output_20)) # (!\ShiftLeft0~89_combout  & ((alu_a_mux_output_22)))))

	.dataa(alu_a_mux_output_20),
	.datab(alu_a_mux_output_22),
	.datac(Mux311),
	.datad(\ShiftLeft0~89_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~90 .lut_mask = 16'hFA0C;
defparam \ShiftLeft0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N22
cycloneive_lcell_comb \ShiftLeft0~91 (
// Equation(s):
// \ShiftLeft0~91_combout  = (Mux291 & (((\ShiftLeft0~77_combout ) # (\ShiftLeft0~78_combout )))) # (!Mux291 & (\ShiftLeft0~90_combout ))

	.dataa(Mux291),
	.datab(\ShiftLeft0~90_combout ),
	.datac(\ShiftLeft0~77_combout ),
	.datad(\ShiftLeft0~78_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~91 .lut_mask = 16'hEEE4;
defparam \ShiftLeft0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N24
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (!\ShiftLeft0~10_combout  & (!\ShiftLeft0~26_combout  & (!Mux281 & \ShiftLeft0~36_combout )))

	.dataa(\ShiftLeft0~10_combout ),
	.datab(\ShiftLeft0~26_combout ),
	.datac(Mux281),
	.datad(\ShiftLeft0~36_combout ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'h0100;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N26
cycloneive_lcell_comb \Mux9~2 (
// Equation(s):
// \Mux9~2_combout  = (\Mux12~2_combout  & (\ShiftRight0~102_combout  & (\Mux12~1_combout ))) # (!\Mux12~2_combout  & (((\Mux9~1_combout ) # (!\Mux12~1_combout ))))

	.dataa(\Mux12~2_combout ),
	.datab(\ShiftRight0~102_combout ),
	.datac(\Mux12~1_combout ),
	.datad(\Mux9~1_combout ),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~2 .lut_mask = 16'hD585;
defparam \Mux9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y41_N2
cycloneive_lcell_comb \Mux9~3 (
// Equation(s):
// \Mux9~3_combout  = (\Mux12~0_combout  & (((\Mux9~2_combout )))) # (!\Mux12~0_combout  & ((\Mux9~2_combout  & (\ShiftLeft0~91_combout )) # (!\Mux9~2_combout  & ((\ShiftLeft0~67_combout )))))

	.dataa(\ShiftLeft0~91_combout ),
	.datab(\Mux12~0_combout ),
	.datac(\ShiftLeft0~67_combout ),
	.datad(\Mux9~2_combout ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~3 .lut_mask = 16'hEE30;
defparam \Mux9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N12
cycloneive_lcell_comb \Mux6~6 (
// Equation(s):
// \Mux6~6_combout  = (\Mux19~1_combout  & (((\Mux19~2_combout )))) # (!\Mux19~1_combout  & ((alu_a_mux_output_25 & (!Mux6 & !\Mux19~2_combout )) # (!alu_a_mux_output_25 & (Mux6 $ (\Mux19~2_combout )))))

	.dataa(alu_a_mux_output_25),
	.datab(Mux6),
	.datac(\Mux19~1_combout ),
	.datad(\Mux19~2_combout ),
	.cin(gnd),
	.combout(\Mux6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~6 .lut_mask = 16'hF106;
defparam \Mux6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N20
cycloneive_lcell_comb \ShiftLeft0~92 (
// Equation(s):
// \ShiftLeft0~92_combout  = (Mux301 & ((alu_a_mux_output_22) # ((!Mux311)))) # (!Mux301 & (((alu_a_mux_output_24 & Mux311))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_22),
	.datac(alu_a_mux_output_24),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftLeft0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~92 .lut_mask = 16'hD8AA;
defparam \ShiftLeft0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N2
cycloneive_lcell_comb \ShiftLeft0~93 (
// Equation(s):
// \ShiftLeft0~93_combout  = (\ShiftLeft0~92_combout  & (((alu_a_mux_output_23) # (Mux311)))) # (!\ShiftLeft0~92_combout  & (alu_a_mux_output_25 & ((!Mux311))))

	.dataa(alu_a_mux_output_25),
	.datab(\ShiftLeft0~92_combout ),
	.datac(alu_a_mux_output_23),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftLeft0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~93 .lut_mask = 16'hCCE2;
defparam \ShiftLeft0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N0
cycloneive_lcell_comb \Mux6~2 (
// Equation(s):
// \Mux6~2_combout  = (\Mux27~2_combout  & (\Mux27~3_combout )) # (!\Mux27~2_combout  & ((\Mux27~3_combout  & (\ShiftLeft0~70_combout )) # (!\Mux27~3_combout  & ((\ShiftLeft0~93_combout )))))

	.dataa(\Mux27~2_combout ),
	.datab(\Mux27~3_combout ),
	.datac(\ShiftLeft0~70_combout ),
	.datad(\ShiftLeft0~93_combout ),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~2 .lut_mask = 16'hD9C8;
defparam \Mux6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N20
cycloneive_lcell_comb \Mux6~3 (
// Equation(s):
// \Mux6~3_combout  = (\Mux27~2_combout  & ((\Mux6~2_combout  & ((\ShiftLeft0~41_combout ))) # (!\Mux6~2_combout  & (\ShiftLeft0~84_combout )))) # (!\Mux27~2_combout  & (((\Mux6~2_combout ))))

	.dataa(\ShiftLeft0~84_combout ),
	.datab(\Mux27~2_combout ),
	.datac(\Mux6~2_combout ),
	.datad(\ShiftLeft0~41_combout ),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~3 .lut_mask = 16'hF838;
defparam \Mux6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N18
cycloneive_lcell_comb \Mux6~8 (
// Equation(s):
// \Mux6~8_combout  = (!\ShiftLeft0~8_combout  & (\Mux6~3_combout  & (!\ShiftLeft0~10_combout  & !\ShiftLeft0~7_combout )))

	.dataa(\ShiftLeft0~8_combout ),
	.datab(\Mux6~3_combout ),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\ShiftLeft0~7_combout ),
	.cin(gnd),
	.combout(\Mux6~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~8 .lut_mask = 16'h0004;
defparam \Mux6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N6
cycloneive_lcell_comb \ShiftRight0~103 (
// Equation(s):
// \ShiftRight0~103_combout  = (!Mux281 & ((Mux291 & (\ShiftRight0~18_combout )) # (!Mux291 & ((\ShiftRight0~20_combout )))))

	.dataa(\ShiftRight0~18_combout ),
	.datab(Mux281),
	.datac(\ShiftRight0~20_combout ),
	.datad(Mux291),
	.cin(gnd),
	.combout(\ShiftRight0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~103 .lut_mask = 16'h2230;
defparam \ShiftRight0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N28
cycloneive_lcell_comb \Mux6~4 (
// Equation(s):
// \Mux6~4_combout  = (\Mux7~0_combout  & ((temp_ALUop_output_0 & ((\ShiftRight0~103_combout ))) # (!temp_ALUop_output_0 & (\Mux6~8_combout )))) # (!\Mux7~0_combout  & (((!temp_ALUop_output_0))))

	.dataa(\Mux7~0_combout ),
	.datab(\Mux6~8_combout ),
	.datac(temp_ALUop_output_0),
	.datad(\ShiftRight0~103_combout ),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~4 .lut_mask = 16'hAD0D;
defparam \Mux6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N26
cycloneive_lcell_comb \Mux6~5 (
// Equation(s):
// \Mux6~5_combout  = (temp_ALUop_output_1 & ((alu_a_mux_output_25 & ((Mux6) # (!\Mux6~4_combout ))) # (!alu_a_mux_output_25 & (Mux6 & !\Mux6~4_combout )))) # (!temp_ALUop_output_1 & (((\Mux6~4_combout ))))

	.dataa(alu_a_mux_output_25),
	.datab(Mux6),
	.datac(temp_ALUop_output_1),
	.datad(\Mux6~4_combout ),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~5 .lut_mask = 16'h8FE0;
defparam \Mux6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N30
cycloneive_lcell_comb \Add0~81 (
// Equation(s):
// \Add0~81_combout  = temp_ALUop_output_0 $ (Mux6)

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(Mux6),
	.cin(gnd),
	.combout(\Add0~81_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~81 .lut_mask = 16'h0FF0;
defparam \Add0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N28
cycloneive_lcell_comb \Add0~82 (
// Equation(s):
// \Add0~82_combout  = temp_ALUop_output_0 $ (Mux7)

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(Mux7),
	.cin(gnd),
	.combout(\Add0~82_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~82 .lut_mask = 16'h0FF0;
defparam \Add0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N2
cycloneive_lcell_comb \Add0~83 (
// Equation(s):
// \Add0~83_combout  = (alu_a_mux_output_24 & ((\Add0~82_combout  & (\Add0~80  & VCC)) # (!\Add0~82_combout  & (!\Add0~80 )))) # (!alu_a_mux_output_24 & ((\Add0~82_combout  & (!\Add0~80 )) # (!\Add0~82_combout  & ((\Add0~80 ) # (GND)))))
// \Add0~84  = CARRY((alu_a_mux_output_24 & (!\Add0~82_combout  & !\Add0~80 )) # (!alu_a_mux_output_24 & ((!\Add0~80 ) # (!\Add0~82_combout ))))

	.dataa(alu_a_mux_output_24),
	.datab(\Add0~82_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~80 ),
	.combout(\Add0~83_combout ),
	.cout(\Add0~84 ));
// synopsys translate_off
defparam \Add0~83 .lut_mask = 16'h9617;
defparam \Add0~83 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N4
cycloneive_lcell_comb \Add0~85 (
// Equation(s):
// \Add0~85_combout  = ((alu_a_mux_output_25 $ (\Add0~81_combout  $ (!\Add0~84 )))) # (GND)
// \Add0~86  = CARRY((alu_a_mux_output_25 & ((\Add0~81_combout ) # (!\Add0~84 ))) # (!alu_a_mux_output_25 & (\Add0~81_combout  & !\Add0~84 )))

	.dataa(alu_a_mux_output_25),
	.datab(\Add0~81_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~84 ),
	.combout(\Add0~85_combout ),
	.cout(\Add0~86 ));
// synopsys translate_off
defparam \Add0~85 .lut_mask = 16'h698E;
defparam \Add0~85 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N24
cycloneive_lcell_comb \ShiftLeft0~50 (
// Equation(s):
// \ShiftLeft0~50_combout  = (Mux281 & (((!Mux291 & \ShiftLeft0~30_combout )))) # (!Mux281 & (\ShiftLeft0~49_combout ))

	.dataa(\ShiftLeft0~49_combout ),
	.datab(Mux291),
	.datac(Mux281),
	.datad(\ShiftLeft0~30_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~50 .lut_mask = 16'h3A0A;
defparam \ShiftLeft0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N4
cycloneive_lcell_comb \Mux4~3 (
// Equation(s):
// \Mux4~3_combout  = (\Mux4~2_combout  & ((\ShiftLeft0~50_combout ) # ((!\Mux27~2_combout )))) # (!\Mux4~2_combout  & (((\Mux27~2_combout  & \ShiftLeft0~87_combout ))))

	.dataa(\Mux4~2_combout ),
	.datab(\ShiftLeft0~50_combout ),
	.datac(\Mux27~2_combout ),
	.datad(\ShiftLeft0~87_combout ),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~3 .lut_mask = 16'hDA8A;
defparam \Mux4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N26
cycloneive_lcell_comb \Mux4~8 (
// Equation(s):
// \Mux4~8_combout  = (!\ShiftLeft0~8_combout  & (!\ShiftLeft0~10_combout  & (\Mux4~3_combout  & !\ShiftLeft0~7_combout )))

	.dataa(\ShiftLeft0~8_combout ),
	.datab(\ShiftLeft0~10_combout ),
	.datac(\Mux4~3_combout ),
	.datad(\ShiftLeft0~7_combout ),
	.cin(gnd),
	.combout(\Mux4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~8 .lut_mask = 16'h0010;
defparam \Mux4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N0
cycloneive_lcell_comb \Mux4~4 (
// Equation(s):
// \Mux4~4_combout  = (\Mux7~0_combout  & ((temp_ALUop_output_0 & ((\ShiftRight0~105_combout ))) # (!temp_ALUop_output_0 & (\Mux4~8_combout )))) # (!\Mux7~0_combout  & (((!temp_ALUop_output_0))))

	.dataa(\Mux7~0_combout ),
	.datab(\Mux4~8_combout ),
	.datac(temp_ALUop_output_0),
	.datad(\ShiftRight0~105_combout ),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~4 .lut_mask = 16'hAD0D;
defparam \Mux4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N6
cycloneive_lcell_comb \Mux4~5 (
// Equation(s):
// \Mux4~5_combout  = (\Mux4~4_combout  & (((Mux4 & alu_a_mux_output_27)) # (!temp_ALUop_output_1))) # (!\Mux4~4_combout  & (temp_ALUop_output_1 & ((Mux4) # (alu_a_mux_output_27))))

	.dataa(\Mux4~4_combout ),
	.datab(temp_ALUop_output_1),
	.datac(Mux4),
	.datad(alu_a_mux_output_27),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~5 .lut_mask = 16'hE662;
defparam \Mux4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N22
cycloneive_lcell_comb \Add0~90 (
// Equation(s):
// \Add0~90_combout  = temp_ALUop_output_0 $ (Mux4)

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(Mux4),
	.cin(gnd),
	.combout(\Add0~90_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~90 .lut_mask = 16'h0FF0;
defparam \Add0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N6
cycloneive_lcell_comb \Add0~88 (
// Equation(s):
// \Add0~88_combout  = (\Add0~87_combout  & ((alu_a_mux_output_26 & (\Add0~86  & VCC)) # (!alu_a_mux_output_26 & (!\Add0~86 )))) # (!\Add0~87_combout  & ((alu_a_mux_output_26 & (!\Add0~86 )) # (!alu_a_mux_output_26 & ((\Add0~86 ) # (GND)))))
// \Add0~89  = CARRY((\Add0~87_combout  & (!alu_a_mux_output_26 & !\Add0~86 )) # (!\Add0~87_combout  & ((!\Add0~86 ) # (!alu_a_mux_output_26))))

	.dataa(\Add0~87_combout ),
	.datab(alu_a_mux_output_26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~86 ),
	.combout(\Add0~88_combout ),
	.cout(\Add0~89 ));
// synopsys translate_off
defparam \Add0~88 .lut_mask = 16'h9617;
defparam \Add0~88 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N8
cycloneive_lcell_comb \Add0~91 (
// Equation(s):
// \Add0~91_combout  = ((\Add0~90_combout  $ (alu_a_mux_output_27 $ (!\Add0~89 )))) # (GND)
// \Add0~92  = CARRY((\Add0~90_combout  & ((alu_a_mux_output_27) # (!\Add0~89 ))) # (!\Add0~90_combout  & (alu_a_mux_output_27 & !\Add0~89 )))

	.dataa(\Add0~90_combout ),
	.datab(alu_a_mux_output_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~89 ),
	.combout(\Add0~91_combout ),
	.cout(\Add0~92 ));
// synopsys translate_off
defparam \Add0~91 .lut_mask = 16'h698E;
defparam \Add0~91 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X68_Y43_N18
cycloneive_lcell_comb \Mux4~6 (
// Equation(s):
// \Mux4~6_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!Mux4 & !alu_a_mux_output_27)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (Mux4 $ (alu_a_mux_output_27))))

	.dataa(\Mux19~2_combout ),
	.datab(Mux4),
	.datac(\Mux19~1_combout ),
	.datad(alu_a_mux_output_27),
	.cin(gnd),
	.combout(\Mux4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~6 .lut_mask = 16'hA1A6;
defparam \Mux4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N18
cycloneive_lcell_comb \ShiftLeft0~102 (
// Equation(s):
// \ShiftLeft0~102_combout  = (Mux311 & (alu_a_mux_output_28)) # (!Mux311 & ((alu_a_mux_output_29)))

	.dataa(gnd),
	.datab(alu_a_mux_output_28),
	.datac(Mux311),
	.datad(alu_a_mux_output_29),
	.cin(gnd),
	.combout(\ShiftLeft0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~102 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N16
cycloneive_lcell_comb \Mux2~3 (
// Equation(s):
// \Mux2~3_combout  = (\ShiftRight0~59_combout  & (\ShiftLeft0~102_combout  & (!\Mux29~0_combout ))) # (!\ShiftRight0~59_combout  & (((\Mux29~0_combout ) # (\ShiftLeft0~93_combout ))))

	.dataa(\ShiftRight0~59_combout ),
	.datab(\ShiftLeft0~102_combout ),
	.datac(\Mux29~0_combout ),
	.datad(\ShiftLeft0~93_combout ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~3 .lut_mask = 16'h5D58;
defparam \Mux2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N2
cycloneive_lcell_comb \Mux2~4 (
// Equation(s):
// \Mux2~4_combout  = (\Mux2~3_combout  & (((\ShiftLeft0~85_combout ) # (!\Mux29~0_combout )))) # (!\Mux2~3_combout  & (\ShiftLeft0~100_combout  & (\Mux29~0_combout )))

	.dataa(\ShiftLeft0~100_combout ),
	.datab(\Mux2~3_combout ),
	.datac(\Mux29~0_combout ),
	.datad(\ShiftLeft0~85_combout ),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~4 .lut_mask = 16'hEC2C;
defparam \Mux2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N24
cycloneive_lcell_comb \Mux2~6 (
// Equation(s):
// \Mux2~6_combout  = (temp_ALUop_output_1) # ((!temp_ALUop_output_0 & Mux271))

	.dataa(temp_ALUop_output_0),
	.datab(temp_ALUop_output_1),
	.datac(gnd),
	.datad(Mux271),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~6 .lut_mask = 16'hDDCC;
defparam \Mux2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N6
cycloneive_lcell_comb \OUTPUT~2 (
// Equation(s):
// \OUTPUT~2_combout  = (Mux2 & alu_a_mux_output_29)

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux2),
	.datad(alu_a_mux_output_29),
	.cin(gnd),
	.combout(\OUTPUT~2_combout ),
	.cout());
// synopsys translate_off
defparam \OUTPUT~2 .lut_mask = 16'hF000;
defparam \OUTPUT~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N2
cycloneive_lcell_comb \Mux2~7 (
// Equation(s):
// \Mux2~7_combout  = (\Mux2~5_combout  & ((\Mux2~6_combout  & (\OUTPUT~2_combout )) # (!\Mux2~6_combout  & ((\ShiftRight0~111_combout ))))) # (!\Mux2~5_combout  & (\Mux2~6_combout ))

	.dataa(\Mux2~5_combout ),
	.datab(\Mux2~6_combout ),
	.datac(\OUTPUT~2_combout ),
	.datad(\ShiftRight0~111_combout ),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~7 .lut_mask = 16'hE6C4;
defparam \Mux2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N22
cycloneive_lcell_comb \Mux2~8 (
// Equation(s):
// \Mux2~8_combout  = (\Mux2~2_combout  & (((\Mux2~7_combout )))) # (!\Mux2~2_combout  & ((\Mux2~7_combout  & (\ShiftLeft0~58_combout )) # (!\Mux2~7_combout  & ((\Mux2~4_combout )))))

	.dataa(\Mux2~2_combout ),
	.datab(\ShiftLeft0~58_combout ),
	.datac(\Mux2~4_combout ),
	.datad(\Mux2~7_combout ),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~8 .lut_mask = 16'hEE50;
defparam \Mux2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N12
cycloneive_lcell_comb \Mux2~9 (
// Equation(s):
// \Mux2~9_combout  = (\Mux2~15_combout  & (!\Mux19~2_combout  & \Mux2~8_combout )) # (!\Mux2~15_combout  & (\Mux19~2_combout ))

	.dataa(\Mux2~15_combout ),
	.datab(gnd),
	.datac(\Mux19~2_combout ),
	.datad(\Mux2~8_combout ),
	.cin(gnd),
	.combout(\Mux2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~9 .lut_mask = 16'h5A50;
defparam \Mux2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N22
cycloneive_lcell_comb \Mux2~10 (
// Equation(s):
// \Mux2~10_combout  = (\Mux19~1_combout  & (((\Mux2~9_combout )))) # (!\Mux19~1_combout  & ((alu_a_mux_output_29 & (!Mux2 & !\Mux2~9_combout )) # (!alu_a_mux_output_29 & (Mux2 $ (\Mux2~9_combout )))))

	.dataa(alu_a_mux_output_29),
	.datab(Mux2),
	.datac(\Mux19~1_combout ),
	.datad(\Mux2~9_combout ),
	.cin(gnd),
	.combout(\Mux2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~10 .lut_mask = 16'hF106;
defparam \Mux2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N16
cycloneive_lcell_comb \Mux2~11 (
// Equation(s):
// \Mux2~11_combout  = (\Mux19~2_combout ) # ((\Mux2~15_combout  & \Mux2~8_combout ))

	.dataa(\Mux2~15_combout ),
	.datab(gnd),
	.datac(\Mux19~2_combout ),
	.datad(\Mux2~8_combout ),
	.cin(gnd),
	.combout(\Mux2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~11 .lut_mask = 16'hFAF0;
defparam \Mux2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N18
cycloneive_lcell_comb \Mux2~12 (
// Equation(s):
// \Mux2~12_combout  = (\Mux19~1_combout  & (((\Mux2~11_combout )))) # (!\Mux19~1_combout  & ((alu_a_mux_output_29 & (!Mux2 & !\Mux2~11_combout )) # (!alu_a_mux_output_29 & (Mux2 $ (\Mux2~11_combout )))))

	.dataa(alu_a_mux_output_29),
	.datab(Mux2),
	.datac(\Mux19~1_combout ),
	.datad(\Mux2~11_combout ),
	.cin(gnd),
	.combout(\Mux2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~12 .lut_mask = 16'hF106;
defparam \Mux2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N4
cycloneive_lcell_comb \Mux2~13 (
// Equation(s):
// \Mux2~13_combout  = (\Mux29~11_combout  & ((alu_a_mux_output_29) # ((Mux2)))) # (!\Mux29~11_combout  & (((\Mux2~12_combout ))))

	.dataa(alu_a_mux_output_29),
	.datab(\Mux2~12_combout ),
	.datac(Mux2),
	.datad(\Mux29~11_combout ),
	.cin(gnd),
	.combout(\Mux2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~13 .lut_mask = 16'hFACC;
defparam \Mux2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N20
cycloneive_lcell_comb \Add0~93 (
// Equation(s):
// \Add0~93_combout  = Mux2 $ (temp_ALUop_output_0)

	.dataa(gnd),
	.datab(Mux2),
	.datac(temp_ALUop_output_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add0~93_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~93 .lut_mask = 16'h3C3C;
defparam \Add0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N10
cycloneive_lcell_comb \Add0~95 (
// Equation(s):
// \Add0~95_combout  = (\Add0~94_combout  & ((alu_a_mux_output_28 & (\Add0~92  & VCC)) # (!alu_a_mux_output_28 & (!\Add0~92 )))) # (!\Add0~94_combout  & ((alu_a_mux_output_28 & (!\Add0~92 )) # (!alu_a_mux_output_28 & ((\Add0~92 ) # (GND)))))
// \Add0~96  = CARRY((\Add0~94_combout  & (!alu_a_mux_output_28 & !\Add0~92 )) # (!\Add0~94_combout  & ((!\Add0~92 ) # (!alu_a_mux_output_28))))

	.dataa(\Add0~94_combout ),
	.datab(alu_a_mux_output_28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~92 ),
	.combout(\Add0~95_combout ),
	.cout(\Add0~96 ));
// synopsys translate_off
defparam \Add0~95 .lut_mask = 16'h9617;
defparam \Add0~95 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N12
cycloneive_lcell_comb \Add0~97 (
// Equation(s):
// \Add0~97_combout  = ((\Add0~93_combout  $ (alu_a_mux_output_29 $ (!\Add0~96 )))) # (GND)
// \Add0~98  = CARRY((\Add0~93_combout  & ((alu_a_mux_output_29) # (!\Add0~96 ))) # (!\Add0~93_combout  & (alu_a_mux_output_29 & !\Add0~96 )))

	.dataa(\Add0~93_combout ),
	.datab(alu_a_mux_output_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~96 ),
	.combout(\Add0~97_combout ),
	.cout(\Add0~98 ));
// synopsys translate_off
defparam \Add0~97 .lut_mask = 16'h698E;
defparam \Add0~97 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N22
cycloneive_lcell_comb \Mux2~5 (
// Equation(s):
// \Mux2~5_combout  = (temp_ALUop_output_1) # ((temp_ALUop_output_0 & \Mux19~0_combout ))

	.dataa(temp_ALUop_output_0),
	.datab(temp_ALUop_output_1),
	.datac(\Mux19~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~5 .lut_mask = 16'hECEC;
defparam \Mux2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N20
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (\Mux2~5_combout  & ((\Mux2~6_combout  & (\OUTPUT~3_combout )) # (!\Mux2~6_combout  & ((\ShiftRight0~108_combout ))))) # (!\Mux2~5_combout  & (((\Mux2~6_combout ))))

	.dataa(\OUTPUT~3_combout ),
	.datab(\ShiftRight0~108_combout ),
	.datac(\Mux2~5_combout ),
	.datad(\Mux2~6_combout ),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hAFC0;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y42_N12
cycloneive_lcell_comb \Mux2~2 (
// Equation(s):
// \Mux2~2_combout  = (temp_ALUop_output_0) # (temp_ALUop_output_1)

	.dataa(gnd),
	.datab(temp_ALUop_output_0),
	.datac(temp_ALUop_output_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~2 .lut_mask = 16'hFCFC;
defparam \Mux2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N24
cycloneive_lcell_comb \ShiftLeft0~61 (
// Equation(s):
// \ShiftLeft0~61_combout  = (Mux281 & ((\ShiftLeft0~29_combout ))) # (!Mux281 & (\ShiftLeft0~60_combout ))

	.dataa(\ShiftLeft0~60_combout ),
	.datab(gnd),
	.datac(Mux281),
	.datad(\ShiftLeft0~29_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~61 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N6
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// \Mux3~3_combout  = (\Mux3~2_combout  & (((\Mux2~2_combout ) # (\ShiftLeft0~61_combout )))) # (!\Mux3~2_combout  & (\Mux3~1_combout  & (!\Mux2~2_combout )))

	.dataa(\Mux3~1_combout ),
	.datab(\Mux3~2_combout ),
	.datac(\Mux2~2_combout ),
	.datad(\ShiftLeft0~61_combout ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hCEC2;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N24
cycloneive_lcell_comb \Mux3~4 (
// Equation(s):
// \Mux3~4_combout  = (\Mux2~15_combout  & (!\Mux19~2_combout  & \Mux3~3_combout )) # (!\Mux2~15_combout  & (\Mux19~2_combout ))

	.dataa(\Mux2~15_combout ),
	.datab(gnd),
	.datac(\Mux19~2_combout ),
	.datad(\Mux3~3_combout ),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~4 .lut_mask = 16'h5A50;
defparam \Mux3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N26
cycloneive_lcell_comb \Mux3~5 (
// Equation(s):
// \Mux3~5_combout  = (\Mux19~1_combout  & (((\Mux3~4_combout )))) # (!\Mux19~1_combout  & ((Mux3 & (!\Mux3~4_combout  & !alu_a_mux_output_28)) # (!Mux3 & (\Mux3~4_combout  $ (alu_a_mux_output_28)))))

	.dataa(\Mux19~1_combout ),
	.datab(Mux3),
	.datac(\Mux3~4_combout ),
	.datad(alu_a_mux_output_28),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~5 .lut_mask = 16'hA1B4;
defparam \Mux3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N8
cycloneive_lcell_comb \Mux3~6 (
// Equation(s):
// \Mux3~6_combout  = (\Mux19~2_combout ) # ((\Mux2~15_combout  & \Mux3~3_combout ))

	.dataa(\Mux2~15_combout ),
	.datab(gnd),
	.datac(\Mux19~2_combout ),
	.datad(\Mux3~3_combout ),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~6 .lut_mask = 16'hFAF0;
defparam \Mux3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N10
cycloneive_lcell_comb \Mux3~7 (
// Equation(s):
// \Mux3~7_combout  = (\Mux19~1_combout  & (((\Mux3~6_combout )))) # (!\Mux19~1_combout  & ((Mux3 & (!\Mux3~6_combout  & !alu_a_mux_output_28)) # (!Mux3 & (\Mux3~6_combout  $ (alu_a_mux_output_28)))))

	.dataa(\Mux19~1_combout ),
	.datab(Mux3),
	.datac(\Mux3~6_combout ),
	.datad(alu_a_mux_output_28),
	.cin(gnd),
	.combout(\Mux3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~7 .lut_mask = 16'hA1B4;
defparam \Mux3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N20
cycloneive_lcell_comb \Mux3~8 (
// Equation(s):
// \Mux3~8_combout  = (\Mux29~11_combout  & (((alu_a_mux_output_28) # (Mux3)))) # (!\Mux29~11_combout  & (\Mux3~7_combout ))

	.dataa(\Mux3~7_combout ),
	.datab(alu_a_mux_output_28),
	.datac(Mux3),
	.datad(\Mux29~11_combout ),
	.cin(gnd),
	.combout(\Mux3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~8 .lut_mask = 16'hFCAA;
defparam \Mux3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N24
cycloneive_lcell_comb \Add0~94 (
// Equation(s):
// \Add0~94_combout  = temp_ALUop_output_0 $ (Mux3)

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(Mux3),
	.cin(gnd),
	.combout(\Add0~94_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~94 .lut_mask = 16'h0FF0;
defparam \Add0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N30
cycloneive_lcell_comb \Add0~99 (
// Equation(s):
// \Add0~99_combout  = temp_ALUop_output_0 $ (Mux0)

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(Mux0),
	.cin(gnd),
	.combout(\Add0~99_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~99 .lut_mask = 16'h0FF0;
defparam \Add0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N14
cycloneive_lcell_comb \Add0~101 (
// Equation(s):
// \Add0~101_combout  = (\Add0~100_combout  & ((alu_a_mux_output_30 & (\Add0~98  & VCC)) # (!alu_a_mux_output_30 & (!\Add0~98 )))) # (!\Add0~100_combout  & ((alu_a_mux_output_30 & (!\Add0~98 )) # (!alu_a_mux_output_30 & ((\Add0~98 ) # (GND)))))
// \Add0~102  = CARRY((\Add0~100_combout  & (!alu_a_mux_output_30 & !\Add0~98 )) # (!\Add0~100_combout  & ((!\Add0~98 ) # (!alu_a_mux_output_30))))

	.dataa(\Add0~100_combout ),
	.datab(alu_a_mux_output_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~98 ),
	.combout(\Add0~101_combout ),
	.cout(\Add0~102 ));
// synopsys translate_off
defparam \Add0~101 .lut_mask = 16'h9617;
defparam \Add0~101 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N16
cycloneive_lcell_comb \Add0~103 (
// Equation(s):
// \Add0~103_combout  = \Add0~99_combout  $ (\Add0~102  $ (!alu_a_mux_output_311))

	.dataa(\Add0~99_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(alu_a_mux_output_311),
	.cin(\Add0~102 ),
	.combout(\Add0~103_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~103 .lut_mask = 16'h5AA5;
defparam \Add0~103 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N14
cycloneive_lcell_comb \ShiftRight0~109 (
// Equation(s):
// \ShiftRight0~109_combout  = (!Mux281 & (!Mux291 & \ShiftRight0~80_combout ))

	.dataa(gnd),
	.datab(Mux281),
	.datac(Mux291),
	.datad(\ShiftRight0~80_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~109_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~109 .lut_mask = 16'h0300;
defparam \ShiftRight0~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N12
cycloneive_lcell_comb \Mux0~3 (
// Equation(s):
// \Mux0~3_combout  = (!\ShiftLeft0~11_combout  & ((Mux281 & (\ShiftLeft0~34_combout )) # (!Mux281 & ((\ShiftLeft0~65_combout )))))

	.dataa(\ShiftLeft0~34_combout ),
	.datab(Mux281),
	.datac(\ShiftLeft0~11_combout ),
	.datad(\ShiftLeft0~65_combout ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~3 .lut_mask = 16'h0B08;
defparam \Mux0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y41_N14
cycloneive_lcell_comb \Mux0~4 (
// Equation(s):
// \Mux0~4_combout  = (\Mux12~1_combout  & ((\Mux12~2_combout  & (\ShiftRight0~109_combout )) # (!\Mux12~2_combout  & ((\Mux0~3_combout ))))) # (!\Mux12~1_combout  & (((!\Mux12~2_combout ))))

	.dataa(\Mux12~1_combout ),
	.datab(\ShiftRight0~109_combout ),
	.datac(\Mux12~2_combout ),
	.datad(\Mux0~3_combout ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~4 .lut_mask = 16'h8F85;
defparam \Mux0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N0
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (Mux291) # ((!Mux301 & Mux311))

	.dataa(Mux301),
	.datab(gnd),
	.datac(Mux291),
	.datad(Mux311),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hF5F0;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N2
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (\ShiftLeft0~13_combout  & (((\ShiftLeft0~102_combout ) # (\Mux1~1_combout )))) # (!\ShiftLeft0~13_combout  & (alu_a_mux_output_311 & ((!\Mux1~1_combout ))))

	.dataa(alu_a_mux_output_311),
	.datab(\ShiftLeft0~13_combout ),
	.datac(\ShiftLeft0~102_combout ),
	.datad(\Mux1~1_combout ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hCCE2;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N12
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (\Mux1~1_combout  & ((\Mux0~1_combout  & (\ShiftLeft0~101_combout )) # (!\Mux0~1_combout  & ((alu_a_mux_output_30))))) # (!\Mux1~1_combout  & (((\Mux0~1_combout ))))

	.dataa(\ShiftLeft0~101_combout ),
	.datab(\Mux1~1_combout ),
	.datac(alu_a_mux_output_30),
	.datad(\Mux0~1_combout ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hBBC0;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N18
cycloneive_lcell_comb \Mux0~5 (
// Equation(s):
// \Mux0~5_combout  = (\Mux12~0_combout  & (((\Mux0~4_combout )))) # (!\Mux12~0_combout  & ((\Mux0~4_combout  & ((\Mux0~2_combout ))) # (!\Mux0~4_combout  & (\ShiftLeft0~88_combout ))))

	.dataa(\Mux12~0_combout ),
	.datab(\ShiftLeft0~88_combout ),
	.datac(\Mux0~4_combout ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~5 .lut_mask = 16'hF4A4;
defparam \Mux0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N26
cycloneive_lcell_comb \Mux0~6 (
// Equation(s):
// \Mux0~6_combout  = (\Mux19~2_combout  & ((\Mux19~1_combout ) # ((!Mux0 & !alu_a_mux_output_311)))) # (!\Mux19~2_combout  & (!\Mux19~1_combout  & (Mux0 $ (alu_a_mux_output_311))))

	.dataa(\Mux19~2_combout ),
	.datab(\Mux19~1_combout ),
	.datac(Mux0),
	.datad(alu_a_mux_output_311),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~6 .lut_mask = 16'h899A;
defparam \Mux0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N30
cycloneive_lcell_comb \Equal0~4 (
// Equation(s):
// \Equal0~4_combout  = (!Mux241 & (!Mux61 & !Mux71))

	.dataa(Mux241),
	.datab(Mux61),
	.datac(gnd),
	.datad(Mux71),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~4 .lut_mask = 16'h0011;
defparam \Equal0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N22
cycloneive_lcell_comb \Equal0~5 (
// Equation(s):
// \Equal0~5_combout  = (temp_ALUop_output_3) # ((!Mux41 & (!Mux51 & \Equal0~4_combout )))

	.dataa(Mux41),
	.datab(temp_ALUop_output_3),
	.datac(Mux51),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~5 .lut_mask = 16'hCDCC;
defparam \Equal0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N4
cycloneive_lcell_comb \Mux9~6 (
// Equation(s):
// \Mux9~6_combout  = (!temp_ALUop_output_3 & ((Mux91) # ((!Mux191 & Mux92))))

	.dataa(temp_ALUop_output_3),
	.datab(Mux191),
	.datac(Mux92),
	.datad(Mux91),
	.cin(gnd),
	.combout(\Mux9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~6 .lut_mask = 16'h5510;
defparam \Mux9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N4
cycloneive_lcell_comb \Mux11~6 (
// Equation(s):
// \Mux11~6_combout  = (temp_ALUop_output_2 & (((Mux112)))) # (!temp_ALUop_output_2 & ((temp_ALUop_output_1 & (Mux111)) # (!temp_ALUop_output_1 & ((Mux112)))))

	.dataa(temp_ALUop_output_2),
	.datab(temp_ALUop_output_1),
	.datac(Mux111),
	.datad(Mux112),
	.cin(gnd),
	.combout(\Mux11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~6 .lut_mask = 16'hFB40;
defparam \Mux11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N26
cycloneive_lcell_comb \Equal0~2 (
// Equation(s):
// \Equal0~2_combout  = (temp_ALUop_output_3) # ((!Mux32 & !\Mux11~6_combout ))

	.dataa(Mux32),
	.datab(temp_ALUop_output_3),
	.datac(gnd),
	.datad(\Mux11~6_combout ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~2 .lut_mask = 16'hCCDD;
defparam \Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N24
cycloneive_lcell_comb \Equal0~3 (
// Equation(s):
// \Equal0~3_combout  = (temp_ALUop_output_3) # ((!Mux261 & (!Mux272 & !Mux251)))

	.dataa(Mux261),
	.datab(temp_ALUop_output_3),
	.datac(Mux272),
	.datad(Mux251),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~3 .lut_mask = 16'hCCCD;
defparam \Equal0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N14
cycloneive_lcell_comb \Equal0~6 (
// Equation(s):
// \Equal0~6_combout  = (\Equal0~5_combout  & (!\Mux9~6_combout  & (\Equal0~2_combout  & \Equal0~3_combout )))

	.dataa(\Equal0~5_combout ),
	.datab(\Mux9~6_combout ),
	.datac(\Equal0~2_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~6 .lut_mask = 16'h2000;
defparam \Equal0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N26
cycloneive_lcell_comb \Equal0~7 (
// Equation(s):
// \Equal0~7_combout  = (Mux172) # ((Mux201) # ((Mux211) # (Mux192)))

	.dataa(Mux172),
	.datab(Mux201),
	.datac(Mux211),
	.datad(Mux192),
	.cin(gnd),
	.combout(\Equal0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~7 .lut_mask = 16'hFFFE;
defparam \Equal0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y43_N22
cycloneive_lcell_comb \Equal0~8 (
// Equation(s):
// \Equal0~8_combout  = (Mux202) # ((Mux173) # ((Mux212) # (Mux193)))

	.dataa(Mux202),
	.datab(Mux173),
	.datac(Mux212),
	.datad(Mux193),
	.cin(gnd),
	.combout(\Equal0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~8 .lut_mask = 16'hFFFE;
defparam \Equal0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N10
cycloneive_lcell_comb \Equal0~9 (
// Equation(s):
// \Equal0~9_combout  = (temp_ALUop_output_2 & (((!\Equal0~8_combout )))) # (!temp_ALUop_output_2 & ((temp_ALUop_output_1 & (!\Equal0~7_combout )) # (!temp_ALUop_output_1 & ((!\Equal0~8_combout )))))

	.dataa(temp_ALUop_output_2),
	.datab(\Equal0~7_combout ),
	.datac(\Equal0~8_combout ),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Equal0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~9 .lut_mask = 16'h1B0F;
defparam \Equal0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N26
cycloneive_lcell_comb \Mux1~8 (
// Equation(s):
// \Mux1~8_combout  = (temp_ALUop_output_1 & ((temp_ALUop_output_2 & ((Mux113))) # (!temp_ALUop_output_2 & (Mux110)))) # (!temp_ALUop_output_1 & (((Mux113))))

	.dataa(Mux110),
	.datab(temp_ALUop_output_1),
	.datac(temp_ALUop_output_2),
	.datad(Mux113),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~8 .lut_mask = 16'hFB08;
defparam \Mux1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N18
cycloneive_lcell_comb \Equal0~10 (
// Equation(s):
// \Equal0~10_combout  = (temp_ALUop_output_3) # ((\Equal0~9_combout  & (!\Mux1~8_combout  & !Mux210)))

	.dataa(temp_ALUop_output_3),
	.datab(\Equal0~9_combout ),
	.datac(\Mux1~8_combout ),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Equal0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~10 .lut_mask = 16'hAAAE;
defparam \Equal0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N2
cycloneive_lcell_comb \Mux23~6 (
// Equation(s):
// \Mux23~6_combout  = (Mux232 & ((temp_ALUop_output_2) # (!temp_ALUop_output_1)))

	.dataa(gnd),
	.datab(temp_ALUop_output_1),
	.datac(temp_ALUop_output_2),
	.datad(Mux232),
	.cin(gnd),
	.combout(\Mux23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~6 .lut_mask = 16'hF300;
defparam \Mux23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N16
cycloneive_lcell_comb \Mux22~6 (
// Equation(s):
// \Mux22~6_combout  = (temp_ALUop_output_1 & ((temp_ALUop_output_2 & (Mux222)) # (!temp_ALUop_output_2 & ((Mux221))))) # (!temp_ALUop_output_1 & (((Mux222))))

	.dataa(temp_ALUop_output_1),
	.datab(temp_ALUop_output_2),
	.datac(Mux222),
	.datad(Mux221),
	.cin(gnd),
	.combout(\Mux22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~6 .lut_mask = 16'hF2D0;
defparam \Mux22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N24
cycloneive_lcell_comb \Mux14~5 (
// Equation(s):
// \Mux14~5_combout  = (temp_ALUop_output_2 & (((Mux142)))) # (!temp_ALUop_output_2 & ((temp_ALUop_output_1 & ((Mux141))) # (!temp_ALUop_output_1 & (Mux142))))

	.dataa(temp_ALUop_output_2),
	.datab(temp_ALUop_output_1),
	.datac(Mux142),
	.datad(Mux141),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~5 .lut_mask = 16'hF4B0;
defparam \Mux14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N30
cycloneive_lcell_comb \Mux16~6 (
// Equation(s):
// \Mux16~6_combout  = (temp_ALUop_output_1 & ((temp_ALUop_output_2 & ((Mux163))) # (!temp_ALUop_output_2 & (Mux162)))) # (!temp_ALUop_output_1 & (((Mux163))))

	.dataa(Mux162),
	.datab(temp_ALUop_output_1),
	.datac(Mux163),
	.datad(temp_ALUop_output_2),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~6 .lut_mask = 16'hF0B8;
defparam \Mux16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N14
cycloneive_lcell_comb \Mux18~6 (
// Equation(s):
// \Mux18~6_combout  = (temp_ALUop_output_1 & ((temp_ALUop_output_2 & ((Mux182))) # (!temp_ALUop_output_2 & (Mux181)))) # (!temp_ALUop_output_1 & (((Mux182))))

	.dataa(temp_ALUop_output_1),
	.datab(Mux181),
	.datac(temp_ALUop_output_2),
	.datad(Mux182),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~6 .lut_mask = 16'hFD08;
defparam \Mux18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N6
cycloneive_lcell_comb \Equal0~11 (
// Equation(s):
// \Equal0~11_combout  = (Mux231) # ((\Mux14~5_combout ) # ((\Mux16~6_combout ) # (\Mux18~6_combout )))

	.dataa(Mux231),
	.datab(\Mux14~5_combout ),
	.datac(\Mux16~6_combout ),
	.datad(\Mux18~6_combout ),
	.cin(gnd),
	.combout(\Equal0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~11 .lut_mask = 16'hFFFE;
defparam \Equal0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N8
cycloneive_lcell_comb \Equal0~12 (
// Equation(s):
// \Equal0~12_combout  = (Mux292) # ((Mux282) # ((\Mux22~6_combout ) # (\Equal0~11_combout )))

	.dataa(Mux292),
	.datab(Mux282),
	.datac(\Mux22~6_combout ),
	.datad(\Equal0~11_combout ),
	.cin(gnd),
	.combout(\Equal0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~12 .lut_mask = 16'hFFFE;
defparam \Equal0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N30
cycloneive_lcell_comb \Equal0~13 (
// Equation(s):
// \Equal0~13_combout  = (!Mux302 & ((temp_ALUop_output_3) # ((!\Mux23~6_combout  & !\Equal0~12_combout ))))

	.dataa(temp_ALUop_output_3),
	.datab(\Mux23~6_combout ),
	.datac(\Equal0~12_combout ),
	.datad(Mux302),
	.cin(gnd),
	.combout(\Equal0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~13 .lut_mask = 16'h00AB;
defparam \Equal0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N16
cycloneive_lcell_comb \Mux13~6 (
// Equation(s):
// \Mux13~6_combout  = (temp_ALUop_output_2 & (Mux132)) # (!temp_ALUop_output_2 & ((temp_ALUop_output_1 & ((Mux131))) # (!temp_ALUop_output_1 & (Mux132))))

	.dataa(Mux132),
	.datab(Mux131),
	.datac(temp_ALUop_output_2),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Mux13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~6 .lut_mask = 16'hACAA;
defparam \Mux13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N8
cycloneive_lcell_comb \Mux8~6 (
// Equation(s):
// \Mux8~6_combout  = (temp_ALUop_output_2 & (((Mux82)))) # (!temp_ALUop_output_2 & ((temp_ALUop_output_1 & (Mux81)) # (!temp_ALUop_output_1 & ((Mux82)))))

	.dataa(Mux81),
	.datab(Mux82),
	.datac(temp_ALUop_output_2),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~6 .lut_mask = 16'hCACC;
defparam \Mux8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N2
cycloneive_lcell_comb \Mux12~9 (
// Equation(s):
// \Mux12~9_combout  = (temp_ALUop_output_1 & ((temp_ALUop_output_2 & ((Mux122))) # (!temp_ALUop_output_2 & (Mux121)))) # (!temp_ALUop_output_1 & (((Mux122))))

	.dataa(Mux121),
	.datab(temp_ALUop_output_1),
	.datac(temp_ALUop_output_2),
	.datad(Mux122),
	.cin(gnd),
	.combout(\Mux12~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~9 .lut_mask = 16'hFB08;
defparam \Mux12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N30
cycloneive_lcell_comb \Equal0~14 (
// Equation(s):
// \Equal0~14_combout  = (\Mux10~6_combout ) # ((\Mux13~6_combout ) # ((\Mux8~6_combout ) # (\Mux12~9_combout )))

	.dataa(\Mux10~6_combout ),
	.datab(\Mux13~6_combout ),
	.datac(\Mux8~6_combout ),
	.datad(\Mux12~9_combout ),
	.cin(gnd),
	.combout(\Equal0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~14 .lut_mask = 16'hFFFE;
defparam \Equal0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N28
cycloneive_lcell_comb \Equal0~17 (
// Equation(s):
// \Equal0~17_combout  = (\Mux0~6_combout ) # ((Mux152) # ((\Mux0~5_combout  & \Mux19~1_combout )))

	.dataa(\Mux0~6_combout ),
	.datab(\Mux0~5_combout ),
	.datac(\Mux19~1_combout ),
	.datad(Mux152),
	.cin(gnd),
	.combout(\Equal0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~17 .lut_mask = 16'hFFEA;
defparam \Equal0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N16
cycloneive_lcell_comb \Equal0~19 (
// Equation(s):
// \Equal0~19_combout  = (temp_ALUop_output_3) # ((temp_ALUop_output_1 & (!\Equal0~18_combout )) # (!temp_ALUop_output_1 & ((!\Equal0~17_combout ))))

	.dataa(\Equal0~18_combout ),
	.datab(temp_ALUop_output_1),
	.datac(temp_ALUop_output_3),
	.datad(\Equal0~17_combout ),
	.cin(gnd),
	.combout(\Equal0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~19 .lut_mask = 16'hF4F7;
defparam \Equal0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N0
cycloneive_lcell_comb \Equal0~23 (
// Equation(s):
// \Equal0~23_combout  = (\Mux0~6_combout  & (((temp_ALUop_output_1)) # (!temp_ALUop_output_2))) # (!\Mux0~6_combout  & (((temp_ALUop_output_2 & !temp_ALUop_output_1)) # (!\Mux0~5_combout )))

	.dataa(\Mux0~6_combout ),
	.datab(temp_ALUop_output_2),
	.datac(\Mux0~5_combout ),
	.datad(temp_ALUop_output_1),
	.cin(gnd),
	.combout(\Equal0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~23 .lut_mask = 16'hAF67;
defparam \Equal0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y43_N30
cycloneive_lcell_comb \Equal0~20 (
// Equation(s):
// \Equal0~20_combout  = (\Equal0~19_combout ) # ((\Equal0~16_combout  & (!\Add0~103_combout  & \Equal0~23_combout )))

	.dataa(\Equal0~16_combout ),
	.datab(\Equal0~19_combout ),
	.datac(\Add0~103_combout ),
	.datad(\Equal0~23_combout ),
	.cin(gnd),
	.combout(\Equal0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~20 .lut_mask = 16'hCECC;
defparam \Equal0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y42_N0
cycloneive_lcell_comb \Equal0~21 (
// Equation(s):
// \Equal0~21_combout  = (\Equal0~13_combout  & (\Equal0~20_combout  & ((temp_ALUop_output_3) # (!\Equal0~14_combout ))))

	.dataa(\Equal0~13_combout ),
	.datab(\Equal0~14_combout ),
	.datac(\Equal0~20_combout ),
	.datad(temp_ALUop_output_3),
	.cin(gnd),
	.combout(\Equal0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~21 .lut_mask = 16'hA020;
defparam \Equal0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N16
cycloneive_lcell_comb \Mux1~3 (
// Equation(s):
// \Mux1~3_combout  = (\ShiftLeft0~13_combout  & ((\ShiftLeft0~103_combout ) # ((\Mux1~1_combout )))) # (!\ShiftLeft0~13_combout  & (((alu_a_mux_output_30 & !\Mux1~1_combout ))))

	.dataa(\ShiftLeft0~103_combout ),
	.datab(\ShiftLeft0~13_combout ),
	.datac(alu_a_mux_output_30),
	.datad(\Mux1~1_combout ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~3 .lut_mask = 16'hCCB8;
defparam \Mux1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N14
cycloneive_lcell_comb \Mux1~4 (
// Equation(s):
// \Mux1~4_combout  = (\Mux1~3_combout  & ((\ShiftLeft0~98_combout ) # ((!\Mux1~1_combout )))) # (!\Mux1~3_combout  & (((alu_a_mux_output_29 & \Mux1~1_combout ))))

	.dataa(\ShiftLeft0~98_combout ),
	.datab(\Mux1~3_combout ),
	.datac(alu_a_mux_output_29),
	.datad(\Mux1~1_combout ),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~4 .lut_mask = 16'hB8CC;
defparam \Mux1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N20
cycloneive_lcell_comb \Mux1~5 (
// Equation(s):
// \Mux1~5_combout  = (!\ShiftLeft0~11_combout  & ((Mux281 & ((\ShiftLeft0~36_combout ))) # (!Mux281 & (\ShiftLeft0~67_combout ))))

	.dataa(Mux281),
	.datab(\ShiftLeft0~11_combout ),
	.datac(\ShiftLeft0~67_combout ),
	.datad(\ShiftLeft0~36_combout ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~5 .lut_mask = 16'h3210;
defparam \Mux1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y42_N14
cycloneive_lcell_comb \Mux1~6 (
// Equation(s):
// \Mux1~6_combout  = (\Mux12~2_combout  & (\ShiftRight0~110_combout  & (\Mux12~1_combout ))) # (!\Mux12~2_combout  & (((\Mux1~5_combout ) # (!\Mux12~1_combout ))))

	.dataa(\ShiftRight0~110_combout ),
	.datab(\Mux12~2_combout ),
	.datac(\Mux12~1_combout ),
	.datad(\Mux1~5_combout ),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~6 .lut_mask = 16'hB383;
defparam \Mux1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y42_N14
cycloneive_lcell_comb \Mux1~7 (
// Equation(s):
// \Mux1~7_combout  = (\Mux12~0_combout  & (((\Mux1~6_combout )))) # (!\Mux12~0_combout  & ((\Mux1~6_combout  & ((\Mux1~4_combout ))) # (!\Mux1~6_combout  & (\ShiftLeft0~91_combout ))))

	.dataa(\ShiftLeft0~91_combout ),
	.datab(\Mux12~0_combout ),
	.datac(\Mux1~4_combout ),
	.datad(\Mux1~6_combout ),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~7 .lut_mask = 16'hFC22;
defparam \Mux1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N20
cycloneive_lcell_comb \Mux1~9 (
// Equation(s):
// \Mux1~9_combout  = (alu_a_mux_output_30 & (!\Mux19~2_combout  & ((\Mux19~1_combout ) # (!Mux1)))) # (!alu_a_mux_output_30 & (\Mux19~2_combout  $ (((\Mux19~1_combout ) # (Mux1)))))

	.dataa(alu_a_mux_output_30),
	.datab(\Mux19~1_combout ),
	.datac(\Mux19~2_combout ),
	.datad(Mux1),
	.cin(gnd),
	.combout(\Mux1~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~9 .lut_mask = 16'h0D1E;
defparam \Mux1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N26
cycloneive_lcell_comb \Add0~100 (
// Equation(s):
// \Add0~100_combout  = Mux1 $ (temp_ALUop_output_0)

	.dataa(Mux1),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add0~100_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~100 .lut_mask = 16'h5A5A;
defparam \Add0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N0
cycloneive_lcell_comb \Mux5~7 (
// Equation(s):
// \Mux5~7_combout  = (\Mux19~2_combout  & (!alu_a_mux_output_26 & (!\Mux19~1_combout  & !Mux5))) # (!\Mux19~2_combout  & ((\Mux19~1_combout ) # (alu_a_mux_output_26 $ (Mux5))))

	.dataa(\Mux19~2_combout ),
	.datab(alu_a_mux_output_26),
	.datac(\Mux19~1_combout ),
	.datad(Mux5),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~7 .lut_mask = 16'h5156;
defparam \Mux5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N12
cycloneive_lcell_comb \ShiftRight0~107 (
// Equation(s):
// \ShiftRight0~107_combout  = (\ShiftRight0~106_combout ) # ((\ShiftRight0~59_combout  & ((\ShiftRight0~65_combout ) # (\ShiftRight0~66_combout ))))

	.dataa(\ShiftRight0~106_combout ),
	.datab(\ShiftRight0~65_combout ),
	.datac(\ShiftRight0~59_combout ),
	.datad(\ShiftRight0~66_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~107_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~107 .lut_mask = 16'hFAEA;
defparam \ShiftRight0~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N8
cycloneive_lcell_comb \ShiftLeft0~96 (
// Equation(s):
// \ShiftLeft0~96_combout  = (Mux301 & ((Mux311 & (alu_a_mux_output_23)) # (!Mux311 & ((alu_a_mux_output_24)))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_23),
	.datac(alu_a_mux_output_24),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftLeft0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~96 .lut_mask = 16'h88A0;
defparam \ShiftLeft0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N10
cycloneive_lcell_comb \ShiftLeft0~97 (
// Equation(s):
// \ShiftLeft0~97_combout  = (Mux311 & ((alu_a_mux_output_25))) # (!Mux311 & (alu_a_mux_output_26))

	.dataa(Mux311),
	.datab(gnd),
	.datac(alu_a_mux_output_26),
	.datad(alu_a_mux_output_25),
	.cin(gnd),
	.combout(\ShiftLeft0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~97 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N4
cycloneive_lcell_comb \ShiftLeft0~98 (
// Equation(s):
// \ShiftLeft0~98_combout  = (\ShiftLeft0~96_combout ) # ((!Mux301 & \ShiftLeft0~97_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~96_combout ),
	.datac(Mux301),
	.datad(\ShiftLeft0~97_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~98 .lut_mask = 16'hCFCC;
defparam \ShiftLeft0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N0
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (\Mux27~2_combout  & ((\ShiftLeft0~90_combout ) # ((\Mux27~3_combout )))) # (!\Mux27~2_combout  & (((\ShiftLeft0~98_combout  & !\Mux27~3_combout ))))

	.dataa(\ShiftLeft0~90_combout ),
	.datab(\Mux27~2_combout ),
	.datac(\ShiftLeft0~98_combout ),
	.datad(\Mux27~3_combout ),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'hCCB8;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N28
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (\Mux5~2_combout  & ((\ShiftLeft0~53_combout ) # ((!\Mux27~3_combout )))) # (!\Mux5~2_combout  & (((\ShiftLeft0~79_combout  & \Mux27~3_combout ))))

	.dataa(\ShiftLeft0~53_combout ),
	.datab(\Mux5~2_combout ),
	.datac(\ShiftLeft0~79_combout ),
	.datad(\Mux27~3_combout ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'hB8CC;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N8
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// \Mux5~6_combout  = (!\ShiftLeft0~8_combout  & (\Mux5~3_combout  & (!\ShiftLeft0~10_combout  & !\ShiftLeft0~7_combout )))

	.dataa(\ShiftLeft0~8_combout ),
	.datab(\Mux5~3_combout ),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\ShiftLeft0~7_combout ),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'h0004;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N2
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (\Mux7~0_combout  & ((temp_ALUop_output_0 & (\ShiftRight0~107_combout )) # (!temp_ALUop_output_0 & ((\Mux5~6_combout ))))) # (!\Mux7~0_combout  & (((!temp_ALUop_output_0))))

	.dataa(\Mux7~0_combout ),
	.datab(\ShiftRight0~107_combout ),
	.datac(temp_ALUop_output_0),
	.datad(\Mux5~6_combout ),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'h8F85;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N8
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (temp_ALUop_output_1 & ((Mux5 & ((alu_a_mux_output_26) # (!\Mux5~4_combout ))) # (!Mux5 & (alu_a_mux_output_26 & !\Mux5~4_combout )))) # (!temp_ALUop_output_1 & (((\Mux5~4_combout ))))

	.dataa(Mux5),
	.datab(alu_a_mux_output_26),
	.datac(temp_ALUop_output_1),
	.datad(\Mux5~4_combout ),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'h8FE0;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N22
cycloneive_lcell_comb \Add0~87 (
// Equation(s):
// \Add0~87_combout  = temp_ALUop_output_0 $ (Mux5)

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_ALUop_output_0),
	.datad(Mux5),
	.cin(gnd),
	.combout(\Add0~87_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~87 .lut_mask = 16'h0FF0;
defparam \Add0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N18
cycloneive_lcell_comb \ShiftRight0~104 (
// Equation(s):
// \ShiftRight0~104_combout  = (!Mux281 & ((Mux291 & ((\ShiftRight0~45_combout ))) # (!Mux291 & (\ShiftRight0~54_combout ))))

	.dataa(\ShiftRight0~54_combout ),
	.datab(\ShiftRight0~45_combout ),
	.datac(Mux281),
	.datad(Mux291),
	.cin(gnd),
	.combout(\ShiftRight0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~104 .lut_mask = 16'h0C0A;
defparam \ShiftRight0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N0
cycloneive_lcell_comb \ShiftLeft0~94 (
// Equation(s):
// \ShiftLeft0~94_combout  = (Mux301 & ((alu_a_mux_output_22) # ((Mux311)))) # (!Mux301 & (((alu_a_mux_output_24 & !Mux311))))

	.dataa(Mux301),
	.datab(alu_a_mux_output_22),
	.datac(alu_a_mux_output_24),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftLeft0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~94 .lut_mask = 16'hAAD8;
defparam \ShiftLeft0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N6
cycloneive_lcell_comb \ShiftLeft0~95 (
// Equation(s):
// \ShiftLeft0~95_combout  = (Mux311 & ((\ShiftLeft0~94_combout  & (alu_a_mux_output_21)) # (!\ShiftLeft0~94_combout  & ((alu_a_mux_output_23))))) # (!Mux311 & (((\ShiftLeft0~94_combout ))))

	.dataa(Mux311),
	.datab(alu_a_mux_output_21),
	.datac(\ShiftLeft0~94_combout ),
	.datad(alu_a_mux_output_23),
	.cin(gnd),
	.combout(\ShiftLeft0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~95 .lut_mask = 16'hDAD0;
defparam \ShiftLeft0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N14
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (\Mux27~2_combout  & (((\ShiftLeft0~81_combout ) # (\Mux27~3_combout )))) # (!\Mux27~2_combout  & (\ShiftLeft0~95_combout  & ((!\Mux27~3_combout ))))

	.dataa(\Mux27~2_combout ),
	.datab(\ShiftLeft0~95_combout ),
	.datac(\ShiftLeft0~81_combout ),
	.datad(\Mux27~3_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hAAE4;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N8
cycloneive_lcell_comb \Mux7~2 (
// Equation(s):
// \Mux7~2_combout  = (\Mux7~1_combout  & (((\ShiftLeft0~45_combout ) # (!\Mux27~3_combout )))) # (!\Mux7~1_combout  & (\ShiftLeft0~73_combout  & ((\Mux27~3_combout ))))

	.dataa(\ShiftLeft0~73_combout ),
	.datab(\ShiftLeft0~45_combout ),
	.datac(\Mux7~1_combout ),
	.datad(\Mux27~3_combout ),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~2 .lut_mask = 16'hCAF0;
defparam \Mux7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N30
cycloneive_lcell_comb \Mux7~3 (
// Equation(s):
// \Mux7~3_combout  = (!\ShiftLeft0~8_combout  & (!\ShiftLeft0~10_combout  & (\Mux7~2_combout  & !\ShiftLeft0~7_combout )))

	.dataa(\ShiftLeft0~8_combout ),
	.datab(\ShiftLeft0~10_combout ),
	.datac(\Mux7~2_combout ),
	.datad(\ShiftLeft0~7_combout ),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~3 .lut_mask = 16'h0010;
defparam \Mux7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N10
cycloneive_lcell_comb \Mux7~4 (
// Equation(s):
// \Mux7~4_combout  = (\Mux7~0_combout  & ((temp_ALUop_output_0 & (\ShiftRight0~104_combout )) # (!temp_ALUop_output_0 & ((\Mux7~3_combout ))))) # (!\Mux7~0_combout  & (((!temp_ALUop_output_0))))

	.dataa(\Mux7~0_combout ),
	.datab(\ShiftRight0~104_combout ),
	.datac(temp_ALUop_output_0),
	.datad(\Mux7~3_combout ),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~4 .lut_mask = 16'h8F85;
defparam \Mux7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N20
cycloneive_lcell_comb \Mux7~5 (
// Equation(s):
// \Mux7~5_combout  = (temp_ALUop_output_1 & ((alu_a_mux_output_24 & ((Mux7) # (!\Mux7~4_combout ))) # (!alu_a_mux_output_24 & (Mux7 & !\Mux7~4_combout )))) # (!temp_ALUop_output_1 & (((\Mux7~4_combout ))))

	.dataa(temp_ALUop_output_1),
	.datab(alu_a_mux_output_24),
	.datac(Mux7),
	.datad(\Mux7~4_combout ),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~5 .lut_mask = 16'hD5A8;
defparam \Mux7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N4
cycloneive_lcell_comb \Mux7~6 (
// Equation(s):
// \Mux7~6_combout  = (\Mux19~2_combout  & (!\Mux19~1_combout  & (!Mux7 & !alu_a_mux_output_24))) # (!\Mux19~2_combout  & ((\Mux19~1_combout ) # (Mux7 $ (alu_a_mux_output_24))))

	.dataa(\Mux19~2_combout ),
	.datab(\Mux19~1_combout ),
	.datac(Mux7),
	.datad(alu_a_mux_output_24),
	.cin(gnd),
	.combout(\Mux7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~6 .lut_mask = 16'h4556;
defparam \Mux7~6 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module alu_a_mux (
	temp_aluResult_1,
	temp_aluResult_0,
	temp_aluResult_2,
	temp_aluResult_3,
	temp_aluResult_5,
	temp_aluResult_4,
	temp_aluResult_7,
	temp_aluResult_6,
	temp_aluResult_9,
	temp_aluResult_8,
	temp_aluResult_11,
	temp_aluResult_10,
	temp_aluResult_13,
	temp_aluResult_12,
	temp_aluResult_15,
	temp_aluResult_14,
	temp_aluResult_17,
	temp_aluResult_16,
	temp_aluResult_19,
	temp_aluResult_18,
	temp_aluResult_20,
	temp_aluResult_21,
	temp_aluResult_23,
	temp_aluResult_22,
	temp_aluResult_25,
	temp_aluResult_24,
	temp_aluResult_26,
	temp_aluResult_27,
	temp_aluResult_29,
	temp_aluResult_28,
	temp_aluResult_31,
	temp_aluResult_30,
	always0,
	Mux30,
	forwarda_1,
	temp_rdat_one_output_1,
	alu_a_mux_output_1,
	Mux31,
	temp_rdat_one_output_0,
	alu_a_mux_output_0,
	Mux29,
	temp_rdat_one_output_2,
	alu_a_mux_output_2,
	Mux27,
	temp_rdat_one_output_4,
	alu_a_mux_output_4,
	Mux28,
	alu_a_mux_output_3,
	temp_rdat_one_output_3,
	alu_a_mux_output_31,
	Mux23,
	temp_rdat_one_output_8,
	alu_a_mux_output_8,
	Mux24,
	temp_rdat_one_output_7,
	alu_a_mux_output_7,
	Mux25,
	temp_rdat_one_output_6,
	alu_a_mux_output_6,
	Mux26,
	temp_rdat_one_output_5,
	alu_a_mux_output_5,
	temp_rdat_one_output_16,
	always01,
	always02,
	Mux15,
	temp_iMemLoad_0,
	alu_a_mux_output_16,
	Mux17,
	temp_rdat_one_output_14,
	alu_a_mux_output_14,
	Mux16,
	temp_rdat_one_output_15,
	alu_a_mux_output_15,
	Mux18,
	temp_rdat_one_output_13,
	alu_a_mux_output_13,
	Mux19,
	temp_rdat_one_output_12,
	alu_a_mux_output_12,
	Mux21,
	temp_rdat_one_output_10,
	alu_a_mux_output_10,
	Mux20,
	temp_rdat_one_output_11,
	alu_a_mux_output_11,
	Mux22,
	temp_rdat_one_output_9,
	alu_a_mux_output_9,
	temp_rdat_one_output_31,
	Mux0,
	temp_iMemLoad_15,
	alu_a_mux_output_311,
	temp_rdat_one_output_30,
	Mux1,
	temp_iMemLoad_14,
	alu_a_mux_output_30,
	temp_rdat_one_output_29,
	Mux2,
	temp_iMemLoad_13,
	alu_a_mux_output_29,
	temp_rdat_one_output_26,
	Mux5,
	temp_iMemLoad_10,
	alu_a_mux_output_26,
	temp_rdat_one_output_25,
	Mux6,
	temp_iMemLoad_9,
	alu_a_mux_output_25,
	temp_rdat_one_output_28,
	Mux3,
	temp_iMemLoad_12,
	alu_a_mux_output_28,
	temp_rdat_one_output_27,
	Mux4,
	temp_iMemLoad_11,
	alu_a_mux_output_27,
	temp_rdat_one_output_17,
	Mux14,
	temp_iMemLoad_1,
	alu_a_mux_output_17,
	temp_rdat_one_output_20,
	Mux11,
	temp_iMemLoad_4,
	alu_a_mux_output_20,
	temp_rdat_one_output_19,
	Mux12,
	temp_iMemLoad_3,
	alu_a_mux_output_19,
	temp_rdat_one_output_18,
	Mux13,
	temp_iMemLoad_2,
	alu_a_mux_output_18,
	temp_rdat_one_output_24,
	Mux7,
	temp_iMemLoad_8,
	alu_a_mux_output_24,
	temp_rdat_one_output_23,
	Mux8,
	temp_iMemLoad_7,
	alu_a_mux_output_23,
	temp_rdat_one_output_22,
	Mux9,
	temp_iMemLoad_6,
	alu_a_mux_output_22,
	temp_rdat_one_output_21,
	Mux10,
	temp_iMemLoad_5,
	alu_a_mux_output_21,
	alu_a_mux_output_32,
	always03,
	devpor,
	devclrn,
	devoe);
input 	temp_aluResult_1;
input 	temp_aluResult_0;
input 	temp_aluResult_2;
input 	temp_aluResult_3;
input 	temp_aluResult_5;
input 	temp_aluResult_4;
input 	temp_aluResult_7;
input 	temp_aluResult_6;
input 	temp_aluResult_9;
input 	temp_aluResult_8;
input 	temp_aluResult_11;
input 	temp_aluResult_10;
input 	temp_aluResult_13;
input 	temp_aluResult_12;
input 	temp_aluResult_15;
input 	temp_aluResult_14;
input 	temp_aluResult_17;
input 	temp_aluResult_16;
input 	temp_aluResult_19;
input 	temp_aluResult_18;
input 	temp_aluResult_20;
input 	temp_aluResult_21;
input 	temp_aluResult_23;
input 	temp_aluResult_22;
input 	temp_aluResult_25;
input 	temp_aluResult_24;
input 	temp_aluResult_26;
input 	temp_aluResult_27;
input 	temp_aluResult_29;
input 	temp_aluResult_28;
input 	temp_aluResult_31;
input 	temp_aluResult_30;
input 	always0;
input 	Mux30;
input 	forwarda_1;
input 	temp_rdat_one_output_1;
output 	alu_a_mux_output_1;
input 	Mux31;
input 	temp_rdat_one_output_0;
output 	alu_a_mux_output_0;
input 	Mux29;
input 	temp_rdat_one_output_2;
output 	alu_a_mux_output_2;
input 	Mux27;
input 	temp_rdat_one_output_4;
output 	alu_a_mux_output_4;
input 	Mux28;
output 	alu_a_mux_output_3;
input 	temp_rdat_one_output_3;
output 	alu_a_mux_output_31;
input 	Mux23;
input 	temp_rdat_one_output_8;
output 	alu_a_mux_output_8;
input 	Mux24;
input 	temp_rdat_one_output_7;
output 	alu_a_mux_output_7;
input 	Mux25;
input 	temp_rdat_one_output_6;
output 	alu_a_mux_output_6;
input 	Mux26;
input 	temp_rdat_one_output_5;
output 	alu_a_mux_output_5;
input 	temp_rdat_one_output_16;
input 	always01;
input 	always02;
input 	Mux15;
input 	temp_iMemLoad_0;
output 	alu_a_mux_output_16;
input 	Mux17;
input 	temp_rdat_one_output_14;
output 	alu_a_mux_output_14;
input 	Mux16;
input 	temp_rdat_one_output_15;
output 	alu_a_mux_output_15;
input 	Mux18;
input 	temp_rdat_one_output_13;
output 	alu_a_mux_output_13;
input 	Mux19;
input 	temp_rdat_one_output_12;
output 	alu_a_mux_output_12;
input 	Mux21;
input 	temp_rdat_one_output_10;
output 	alu_a_mux_output_10;
input 	Mux20;
input 	temp_rdat_one_output_11;
output 	alu_a_mux_output_11;
input 	Mux22;
input 	temp_rdat_one_output_9;
output 	alu_a_mux_output_9;
input 	temp_rdat_one_output_31;
input 	Mux0;
input 	temp_iMemLoad_15;
output 	alu_a_mux_output_311;
input 	temp_rdat_one_output_30;
input 	Mux1;
input 	temp_iMemLoad_14;
output 	alu_a_mux_output_30;
input 	temp_rdat_one_output_29;
input 	Mux2;
input 	temp_iMemLoad_13;
output 	alu_a_mux_output_29;
input 	temp_rdat_one_output_26;
input 	Mux5;
input 	temp_iMemLoad_10;
output 	alu_a_mux_output_26;
input 	temp_rdat_one_output_25;
input 	Mux6;
input 	temp_iMemLoad_9;
output 	alu_a_mux_output_25;
input 	temp_rdat_one_output_28;
input 	Mux3;
input 	temp_iMemLoad_12;
output 	alu_a_mux_output_28;
input 	temp_rdat_one_output_27;
input 	Mux4;
input 	temp_iMemLoad_11;
output 	alu_a_mux_output_27;
input 	temp_rdat_one_output_17;
input 	Mux14;
input 	temp_iMemLoad_1;
output 	alu_a_mux_output_17;
input 	temp_rdat_one_output_20;
input 	Mux11;
input 	temp_iMemLoad_4;
output 	alu_a_mux_output_20;
input 	temp_rdat_one_output_19;
input 	Mux12;
input 	temp_iMemLoad_3;
output 	alu_a_mux_output_19;
input 	temp_rdat_one_output_18;
input 	Mux13;
input 	temp_iMemLoad_2;
output 	alu_a_mux_output_18;
input 	temp_rdat_one_output_24;
input 	Mux7;
input 	temp_iMemLoad_8;
output 	alu_a_mux_output_24;
input 	temp_rdat_one_output_23;
input 	Mux8;
input 	temp_iMemLoad_7;
output 	alu_a_mux_output_23;
input 	temp_rdat_one_output_22;
input 	Mux9;
input 	temp_iMemLoad_6;
output 	alu_a_mux_output_22;
input 	temp_rdat_one_output_21;
input 	Mux10;
input 	temp_iMemLoad_5;
output 	alu_a_mux_output_21;
output 	alu_a_mux_output_32;
input 	always03;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \alu_a_mux_output[1]~0_combout ;
wire \alu_a_mux_output[0]~2_combout ;
wire \alu_a_mux_output[2]~4_combout ;
wire \alu_a_mux_output[4]~6_combout ;
wire \alu_a_mux_output[8]~10_combout ;
wire \alu_a_mux_output[7]~12_combout ;
wire \alu_a_mux_output[6]~14_combout ;
wire \alu_a_mux_output[5]~16_combout ;
wire \alu_a_mux_output[16]~18_combout ;
wire \alu_a_mux_output[16]~19_combout ;
wire \alu_a_mux_output[14]~21_combout ;
wire \alu_a_mux_output[15]~23_combout ;
wire \alu_a_mux_output[13]~25_combout ;
wire \alu_a_mux_output[12]~27_combout ;
wire \alu_a_mux_output[10]~29_combout ;
wire \alu_a_mux_output[11]~31_combout ;
wire \alu_a_mux_output[9]~33_combout ;
wire \alu_a_mux_output[31]~35_combout ;
wire \alu_a_mux_output[30]~37_combout ;
wire \alu_a_mux_output[29]~39_combout ;
wire \alu_a_mux_output[26]~41_combout ;
wire \alu_a_mux_output[25]~43_combout ;
wire \alu_a_mux_output[28]~45_combout ;
wire \alu_a_mux_output[27]~47_combout ;
wire \alu_a_mux_output[17]~49_combout ;
wire \alu_a_mux_output[20]~51_combout ;
wire \alu_a_mux_output[19]~53_combout ;
wire \alu_a_mux_output[18]~55_combout ;
wire \alu_a_mux_output[24]~57_combout ;
wire \alu_a_mux_output[23]~59_combout ;
wire \alu_a_mux_output[22]~61_combout ;
wire \alu_a_mux_output[21]~63_combout ;


// Location: LCCOMB_X66_Y44_N14
cycloneive_lcell_comb \alu_a_mux_output[1]~1 (
// Equation(s):
// alu_a_mux_output_1 = (forwarda_1 & (!always07 & (Mux30))) # (!forwarda_1 & (((\alu_a_mux_output[1]~0_combout ))))

	.dataa(always03),
	.datab(Mux30),
	.datac(forwarda_1),
	.datad(\alu_a_mux_output[1]~0_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_1),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[1]~1 .lut_mask = 16'h4F40;
defparam \alu_a_mux_output[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N0
cycloneive_lcell_comb \alu_a_mux_output[0]~3 (
// Equation(s):
// alu_a_mux_output_0 = (forwarda_1 & (((Mux31 & !always07)))) # (!forwarda_1 & (\alu_a_mux_output[0]~2_combout ))

	.dataa(\alu_a_mux_output[0]~2_combout ),
	.datab(forwarda_1),
	.datac(Mux31),
	.datad(always03),
	.cin(gnd),
	.combout(alu_a_mux_output_0),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[0]~3 .lut_mask = 16'h22E2;
defparam \alu_a_mux_output[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N26
cycloneive_lcell_comb \alu_a_mux_output[2]~5 (
// Equation(s):
// alu_a_mux_output_2 = (forwarda_1 & (Mux29 & ((!always07)))) # (!forwarda_1 & (((\alu_a_mux_output[2]~4_combout ))))

	.dataa(Mux29),
	.datab(\alu_a_mux_output[2]~4_combout ),
	.datac(forwarda_1),
	.datad(always03),
	.cin(gnd),
	.combout(alu_a_mux_output_2),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[2]~5 .lut_mask = 16'h0CAC;
defparam \alu_a_mux_output[2]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N4
cycloneive_lcell_comb \alu_a_mux_output[4]~7 (
// Equation(s):
// alu_a_mux_output_4 = (forwarda_1 & (((Mux27 & !always07)))) # (!forwarda_1 & (\alu_a_mux_output[4]~6_combout ))

	.dataa(\alu_a_mux_output[4]~6_combout ),
	.datab(forwarda_1),
	.datac(Mux27),
	.datad(always03),
	.cin(gnd),
	.combout(alu_a_mux_output_4),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[4]~7 .lut_mask = 16'h22E2;
defparam \alu_a_mux_output[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N0
cycloneive_lcell_comb \alu_a_mux_output[3]~8 (
// Equation(s):
// alu_a_mux_output_3 = (always07 & (temp_aluResult_3 & ((!forwarda_1)))) # (!always07 & (((Mux28 & forwarda_1))))

	.dataa(always03),
	.datab(temp_aluResult_3),
	.datac(Mux28),
	.datad(forwarda_1),
	.cin(gnd),
	.combout(alu_a_mux_output_3),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[3]~8 .lut_mask = 16'h5088;
defparam \alu_a_mux_output[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N28
cycloneive_lcell_comb \alu_a_mux_output[3]~9 (
// Equation(s):
// alu_a_mux_output_31 = (alu_a_mux_output_3) # ((!forwarda_1 & (!always07 & temp_rdat_one_output_3)))

	.dataa(forwarda_1),
	.datab(alu_a_mux_output_3),
	.datac(always03),
	.datad(temp_rdat_one_output_3),
	.cin(gnd),
	.combout(alu_a_mux_output_31),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[3]~9 .lut_mask = 16'hCDCC;
defparam \alu_a_mux_output[3]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N2
cycloneive_lcell_comb \alu_a_mux_output[8]~11 (
// Equation(s):
// alu_a_mux_output_8 = (\alu_a_mux_output[8]~10_combout ) # ((!always07 & (!forwarda_1 & temp_rdat_one_output_8)))

	.dataa(always03),
	.datab(forwarda_1),
	.datac(temp_rdat_one_output_8),
	.datad(\alu_a_mux_output[8]~10_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_8),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[8]~11 .lut_mask = 16'hFF10;
defparam \alu_a_mux_output[8]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N30
cycloneive_lcell_comb \alu_a_mux_output[7]~13 (
// Equation(s):
// alu_a_mux_output_7 = (\alu_a_mux_output[7]~12_combout ) # ((!always07 & (temp_rdat_one_output_7 & !forwarda_1)))

	.dataa(always03),
	.datab(temp_rdat_one_output_7),
	.datac(forwarda_1),
	.datad(\alu_a_mux_output[7]~12_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_7),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[7]~13 .lut_mask = 16'hFF04;
defparam \alu_a_mux_output[7]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N8
cycloneive_lcell_comb \alu_a_mux_output[6]~15 (
// Equation(s):
// alu_a_mux_output_6 = (\alu_a_mux_output[6]~14_combout ) # ((temp_rdat_one_output_6 & (!always07 & !forwarda_1)))

	.dataa(temp_rdat_one_output_6),
	.datab(\alu_a_mux_output[6]~14_combout ),
	.datac(always03),
	.datad(forwarda_1),
	.cin(gnd),
	.combout(alu_a_mux_output_6),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[6]~15 .lut_mask = 16'hCCCE;
defparam \alu_a_mux_output[6]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N0
cycloneive_lcell_comb \alu_a_mux_output[5]~17 (
// Equation(s):
// alu_a_mux_output_5 = (\alu_a_mux_output[5]~16_combout ) # ((!always07 & (!forwarda_1 & temp_rdat_one_output_5)))

	.dataa(always03),
	.datab(forwarda_1),
	.datac(temp_rdat_one_output_5),
	.datad(\alu_a_mux_output[5]~16_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_5),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[5]~17 .lut_mask = 16'hFF10;
defparam \alu_a_mux_output[5]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N16
cycloneive_lcell_comb \alu_a_mux_output[16]~20 (
// Equation(s):
// alu_a_mux_output_16 = (\alu_a_mux_output[16]~18_combout  & ((\alu_a_mux_output[16]~19_combout  & (temp_iMemLoad_0)) # (!\alu_a_mux_output[16]~19_combout  & ((temp_rdat_one_output_16))))) # (!\alu_a_mux_output[16]~18_combout  & 
// (((\alu_a_mux_output[16]~19_combout ))))

	.dataa(temp_iMemLoad_0),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(temp_rdat_one_output_16),
	.datad(\alu_a_mux_output[16]~19_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_16),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[16]~20 .lut_mask = 16'hBBC0;
defparam \alu_a_mux_output[16]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N6
cycloneive_lcell_comb \alu_a_mux_output[14]~22 (
// Equation(s):
// alu_a_mux_output_14 = (\alu_a_mux_output[14]~21_combout ) # ((!forwarda_1 & (temp_rdat_one_output_14 & !always07)))

	.dataa(forwarda_1),
	.datab(temp_rdat_one_output_14),
	.datac(\alu_a_mux_output[14]~21_combout ),
	.datad(always03),
	.cin(gnd),
	.combout(alu_a_mux_output_14),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[14]~22 .lut_mask = 16'hF0F4;
defparam \alu_a_mux_output[14]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N20
cycloneive_lcell_comb \alu_a_mux_output[15]~24 (
// Equation(s):
// alu_a_mux_output_15 = (\alu_a_mux_output[15]~23_combout ) # ((!always07 & (!forwarda_1 & temp_rdat_one_output_15)))

	.dataa(always03),
	.datab(forwarda_1),
	.datac(temp_rdat_one_output_15),
	.datad(\alu_a_mux_output[15]~23_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_15),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[15]~24 .lut_mask = 16'hFF10;
defparam \alu_a_mux_output[15]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N6
cycloneive_lcell_comb \alu_a_mux_output[13]~26 (
// Equation(s):
// alu_a_mux_output_13 = (\alu_a_mux_output[13]~25_combout ) # ((!always07 & (temp_rdat_one_output_13 & !forwarda_1)))

	.dataa(always03),
	.datab(temp_rdat_one_output_13),
	.datac(\alu_a_mux_output[13]~25_combout ),
	.datad(forwarda_1),
	.cin(gnd),
	.combout(alu_a_mux_output_13),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[13]~26 .lut_mask = 16'hF0F4;
defparam \alu_a_mux_output[13]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N10
cycloneive_lcell_comb \alu_a_mux_output[12]~28 (
// Equation(s):
// alu_a_mux_output_12 = (\alu_a_mux_output[12]~27_combout ) # ((!always07 & (!forwarda_1 & temp_rdat_one_output_12)))

	.dataa(\alu_a_mux_output[12]~27_combout ),
	.datab(always03),
	.datac(forwarda_1),
	.datad(temp_rdat_one_output_12),
	.cin(gnd),
	.combout(alu_a_mux_output_12),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[12]~28 .lut_mask = 16'hABAA;
defparam \alu_a_mux_output[12]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N0
cycloneive_lcell_comb \alu_a_mux_output[10]~30 (
// Equation(s):
// alu_a_mux_output_10 = (\alu_a_mux_output[10]~29_combout ) # ((!forwarda_1 & (temp_rdat_one_output_10 & !always07)))

	.dataa(\alu_a_mux_output[10]~29_combout ),
	.datab(forwarda_1),
	.datac(temp_rdat_one_output_10),
	.datad(always03),
	.cin(gnd),
	.combout(alu_a_mux_output_10),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[10]~30 .lut_mask = 16'hAABA;
defparam \alu_a_mux_output[10]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N16
cycloneive_lcell_comb \alu_a_mux_output[11]~32 (
// Equation(s):
// alu_a_mux_output_11 = (\alu_a_mux_output[11]~31_combout ) # ((!forwarda_1 & (temp_rdat_one_output_11 & !always07)))

	.dataa(forwarda_1),
	.datab(temp_rdat_one_output_11),
	.datac(always03),
	.datad(\alu_a_mux_output[11]~31_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_11),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[11]~32 .lut_mask = 16'hFF04;
defparam \alu_a_mux_output[11]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N24
cycloneive_lcell_comb \alu_a_mux_output[9]~34 (
// Equation(s):
// alu_a_mux_output_9 = (\alu_a_mux_output[9]~33_combout ) # ((!always07 & (temp_rdat_one_output_9 & !forwarda_1)))

	.dataa(always03),
	.datab(temp_rdat_one_output_9),
	.datac(\alu_a_mux_output[9]~33_combout ),
	.datad(forwarda_1),
	.cin(gnd),
	.combout(alu_a_mux_output_9),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[9]~34 .lut_mask = 16'hF0F4;
defparam \alu_a_mux_output[9]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N30
cycloneive_lcell_comb \alu_a_mux_output[31]~36 (
// Equation(s):
// alu_a_mux_output_311 = (\alu_a_mux_output[16]~18_combout  & ((\alu_a_mux_output[31]~35_combout  & (temp_iMemLoad_15)) # (!\alu_a_mux_output[31]~35_combout  & ((temp_rdat_one_output_31))))) # (!\alu_a_mux_output[16]~18_combout  & 
// (((\alu_a_mux_output[31]~35_combout ))))

	.dataa(\alu_a_mux_output[16]~18_combout ),
	.datab(temp_iMemLoad_15),
	.datac(\alu_a_mux_output[31]~35_combout ),
	.datad(temp_rdat_one_output_31),
	.cin(gnd),
	.combout(alu_a_mux_output_311),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[31]~36 .lut_mask = 16'hDAD0;
defparam \alu_a_mux_output[31]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N10
cycloneive_lcell_comb \alu_a_mux_output[30]~38 (
// Equation(s):
// alu_a_mux_output_30 = (\alu_a_mux_output[30]~37_combout  & ((temp_iMemLoad_14) # ((!\alu_a_mux_output[16]~18_combout )))) # (!\alu_a_mux_output[30]~37_combout  & (((\alu_a_mux_output[16]~18_combout  & temp_rdat_one_output_30))))

	.dataa(temp_iMemLoad_14),
	.datab(\alu_a_mux_output[30]~37_combout ),
	.datac(\alu_a_mux_output[16]~18_combout ),
	.datad(temp_rdat_one_output_30),
	.cin(gnd),
	.combout(alu_a_mux_output_30),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[30]~38 .lut_mask = 16'hBC8C;
defparam \alu_a_mux_output[30]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N22
cycloneive_lcell_comb \alu_a_mux_output[29]~40 (
// Equation(s):
// alu_a_mux_output_29 = (\alu_a_mux_output[29]~39_combout  & (((temp_iMemLoad_13)) # (!\alu_a_mux_output[16]~18_combout ))) # (!\alu_a_mux_output[29]~39_combout  & (\alu_a_mux_output[16]~18_combout  & ((temp_rdat_one_output_29))))

	.dataa(\alu_a_mux_output[29]~39_combout ),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(temp_iMemLoad_13),
	.datad(temp_rdat_one_output_29),
	.cin(gnd),
	.combout(alu_a_mux_output_29),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[29]~40 .lut_mask = 16'hE6A2;
defparam \alu_a_mux_output[29]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N14
cycloneive_lcell_comb \alu_a_mux_output[26]~42 (
// Equation(s):
// alu_a_mux_output_26 = (\alu_a_mux_output[16]~18_combout  & ((\alu_a_mux_output[26]~41_combout  & (temp_iMemLoad_10)) # (!\alu_a_mux_output[26]~41_combout  & ((temp_rdat_one_output_26))))) # (!\alu_a_mux_output[16]~18_combout  & 
// (((\alu_a_mux_output[26]~41_combout ))))

	.dataa(temp_iMemLoad_10),
	.datab(temp_rdat_one_output_26),
	.datac(\alu_a_mux_output[16]~18_combout ),
	.datad(\alu_a_mux_output[26]~41_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_26),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[26]~42 .lut_mask = 16'hAFC0;
defparam \alu_a_mux_output[26]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N8
cycloneive_lcell_comb \alu_a_mux_output[25]~44 (
// Equation(s):
// alu_a_mux_output_25 = (\alu_a_mux_output[25]~43_combout  & ((temp_iMemLoad_9) # ((!\alu_a_mux_output[16]~18_combout )))) # (!\alu_a_mux_output[25]~43_combout  & (((\alu_a_mux_output[16]~18_combout  & temp_rdat_one_output_25))))

	.dataa(\alu_a_mux_output[25]~43_combout ),
	.datab(temp_iMemLoad_9),
	.datac(\alu_a_mux_output[16]~18_combout ),
	.datad(temp_rdat_one_output_25),
	.cin(gnd),
	.combout(alu_a_mux_output_25),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[25]~44 .lut_mask = 16'hDA8A;
defparam \alu_a_mux_output[25]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N28
cycloneive_lcell_comb \alu_a_mux_output[28]~46 (
// Equation(s):
// alu_a_mux_output_28 = (\alu_a_mux_output[16]~18_combout  & ((\alu_a_mux_output[28]~45_combout  & ((temp_iMemLoad_12))) # (!\alu_a_mux_output[28]~45_combout  & (temp_rdat_one_output_28)))) # (!\alu_a_mux_output[16]~18_combout  & 
// (((\alu_a_mux_output[28]~45_combout ))))

	.dataa(temp_rdat_one_output_28),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(\alu_a_mux_output[28]~45_combout ),
	.datad(temp_iMemLoad_12),
	.cin(gnd),
	.combout(alu_a_mux_output_28),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[28]~46 .lut_mask = 16'hF838;
defparam \alu_a_mux_output[28]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N8
cycloneive_lcell_comb \alu_a_mux_output[27]~48 (
// Equation(s):
// alu_a_mux_output_27 = (\alu_a_mux_output[27]~47_combout  & ((temp_iMemLoad_11) # ((!\alu_a_mux_output[16]~18_combout )))) # (!\alu_a_mux_output[27]~47_combout  & (((\alu_a_mux_output[16]~18_combout  & temp_rdat_one_output_27))))

	.dataa(\alu_a_mux_output[27]~47_combout ),
	.datab(temp_iMemLoad_11),
	.datac(\alu_a_mux_output[16]~18_combout ),
	.datad(temp_rdat_one_output_27),
	.cin(gnd),
	.combout(alu_a_mux_output_27),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[27]~48 .lut_mask = 16'hDA8A;
defparam \alu_a_mux_output[27]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N20
cycloneive_lcell_comb \alu_a_mux_output[17]~50 (
// Equation(s):
// alu_a_mux_output_17 = (\alu_a_mux_output[17]~49_combout  & ((temp_iMemLoad_1) # ((!\alu_a_mux_output[16]~18_combout )))) # (!\alu_a_mux_output[17]~49_combout  & (((temp_rdat_one_output_17 & \alu_a_mux_output[16]~18_combout ))))

	.dataa(temp_iMemLoad_1),
	.datab(temp_rdat_one_output_17),
	.datac(\alu_a_mux_output[17]~49_combout ),
	.datad(\alu_a_mux_output[16]~18_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_17),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[17]~50 .lut_mask = 16'hACF0;
defparam \alu_a_mux_output[17]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N4
cycloneive_lcell_comb \alu_a_mux_output[20]~52 (
// Equation(s):
// alu_a_mux_output_20 = (\alu_a_mux_output[20]~51_combout  & (((temp_iMemLoad_4) # (!\alu_a_mux_output[16]~18_combout )))) # (!\alu_a_mux_output[20]~51_combout  & (temp_rdat_one_output_20 & ((\alu_a_mux_output[16]~18_combout ))))

	.dataa(temp_rdat_one_output_20),
	.datab(\alu_a_mux_output[20]~51_combout ),
	.datac(temp_iMemLoad_4),
	.datad(\alu_a_mux_output[16]~18_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_20),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[20]~52 .lut_mask = 16'hE2CC;
defparam \alu_a_mux_output[20]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N18
cycloneive_lcell_comb \alu_a_mux_output[19]~54 (
// Equation(s):
// alu_a_mux_output_19 = (\alu_a_mux_output[16]~18_combout  & ((\alu_a_mux_output[19]~53_combout  & (temp_iMemLoad_3)) # (!\alu_a_mux_output[19]~53_combout  & ((temp_rdat_one_output_19))))) # (!\alu_a_mux_output[16]~18_combout  & 
// (((\alu_a_mux_output[19]~53_combout ))))

	.dataa(temp_iMemLoad_3),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(temp_rdat_one_output_19),
	.datad(\alu_a_mux_output[19]~53_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_19),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[19]~54 .lut_mask = 16'hBBC0;
defparam \alu_a_mux_output[19]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N6
cycloneive_lcell_comb \alu_a_mux_output[18]~56 (
// Equation(s):
// alu_a_mux_output_18 = (\alu_a_mux_output[16]~18_combout  & ((\alu_a_mux_output[18]~55_combout  & (temp_iMemLoad_2)) # (!\alu_a_mux_output[18]~55_combout  & ((temp_rdat_one_output_18))))) # (!\alu_a_mux_output[16]~18_combout  & 
// (((\alu_a_mux_output[18]~55_combout ))))

	.dataa(temp_iMemLoad_2),
	.datab(temp_rdat_one_output_18),
	.datac(\alu_a_mux_output[16]~18_combout ),
	.datad(\alu_a_mux_output[18]~55_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_18),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[18]~56 .lut_mask = 16'hAFC0;
defparam \alu_a_mux_output[18]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N30
cycloneive_lcell_comb \alu_a_mux_output[24]~58 (
// Equation(s):
// alu_a_mux_output_24 = (\alu_a_mux_output[24]~57_combout  & (((temp_iMemLoad_8)) # (!\alu_a_mux_output[16]~18_combout ))) # (!\alu_a_mux_output[24]~57_combout  & (\alu_a_mux_output[16]~18_combout  & ((temp_rdat_one_output_24))))

	.dataa(\alu_a_mux_output[24]~57_combout ),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(temp_iMemLoad_8),
	.datad(temp_rdat_one_output_24),
	.cin(gnd),
	.combout(alu_a_mux_output_24),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[24]~58 .lut_mask = 16'hE6A2;
defparam \alu_a_mux_output[24]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N8
cycloneive_lcell_comb \alu_a_mux_output[23]~60 (
// Equation(s):
// alu_a_mux_output_23 = (\alu_a_mux_output[23]~59_combout  & (((temp_iMemLoad_7) # (!\alu_a_mux_output[16]~18_combout )))) # (!\alu_a_mux_output[23]~59_combout  & (temp_rdat_one_output_23 & (\alu_a_mux_output[16]~18_combout )))

	.dataa(temp_rdat_one_output_23),
	.datab(\alu_a_mux_output[23]~59_combout ),
	.datac(\alu_a_mux_output[16]~18_combout ),
	.datad(temp_iMemLoad_7),
	.cin(gnd),
	.combout(alu_a_mux_output_23),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[23]~60 .lut_mask = 16'hEC2C;
defparam \alu_a_mux_output[23]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N30
cycloneive_lcell_comb \alu_a_mux_output[22]~62 (
// Equation(s):
// alu_a_mux_output_22 = (\alu_a_mux_output[16]~18_combout  & ((\alu_a_mux_output[22]~61_combout  & (temp_iMemLoad_6)) # (!\alu_a_mux_output[22]~61_combout  & ((temp_rdat_one_output_22))))) # (!\alu_a_mux_output[16]~18_combout  & 
// (((\alu_a_mux_output[22]~61_combout ))))

	.dataa(temp_iMemLoad_6),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(temp_rdat_one_output_22),
	.datad(\alu_a_mux_output[22]~61_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_22),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[22]~62 .lut_mask = 16'hBBC0;
defparam \alu_a_mux_output[22]~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N8
cycloneive_lcell_comb \alu_a_mux_output[21]~64 (
// Equation(s):
// alu_a_mux_output_21 = (\alu_a_mux_output[21]~63_combout  & ((temp_iMemLoad_5) # ((!\alu_a_mux_output[16]~18_combout )))) # (!\alu_a_mux_output[21]~63_combout  & (((temp_rdat_one_output_21 & \alu_a_mux_output[16]~18_combout ))))

	.dataa(temp_iMemLoad_5),
	.datab(\alu_a_mux_output[21]~63_combout ),
	.datac(temp_rdat_one_output_21),
	.datad(\alu_a_mux_output[16]~18_combout ),
	.cin(gnd),
	.combout(alu_a_mux_output_21),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[21]~64 .lut_mask = 16'hB8CC;
defparam \alu_a_mux_output[21]~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N26
cycloneive_lcell_comb \alu_a_mux_output[3]~65 (
// Equation(s):
// alu_a_mux_output_32 = (!forwarda_1 & (temp_rdat_one_output_3 & !always07))

	.dataa(forwarda_1),
	.datab(temp_rdat_one_output_3),
	.datac(always03),
	.datad(gnd),
	.cin(gnd),
	.combout(alu_a_mux_output_32),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[3]~65 .lut_mask = 16'h0404;
defparam \alu_a_mux_output[3]~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N16
cycloneive_lcell_comb \alu_a_mux_output[1]~0 (
// Equation(s):
// \alu_a_mux_output[1]~0_combout  = (always07 & ((temp_aluResult_1))) # (!always07 & (temp_rdat_one_output_1))

	.dataa(temp_rdat_one_output_1),
	.datab(gnd),
	.datac(temp_aluResult_1),
	.datad(always03),
	.cin(gnd),
	.combout(\alu_a_mux_output[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[1]~0 .lut_mask = 16'hF0AA;
defparam \alu_a_mux_output[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N10
cycloneive_lcell_comb \alu_a_mux_output[0]~2 (
// Equation(s):
// \alu_a_mux_output[0]~2_combout  = (always07 & ((temp_aluResult_0))) # (!always07 & (temp_rdat_one_output_0))

	.dataa(gnd),
	.datab(temp_rdat_one_output_0),
	.datac(temp_aluResult_0),
	.datad(always03),
	.cin(gnd),
	.combout(\alu_a_mux_output[0]~2_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[0]~2 .lut_mask = 16'hF0CC;
defparam \alu_a_mux_output[0]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N24
cycloneive_lcell_comb \alu_a_mux_output[2]~4 (
// Equation(s):
// \alu_a_mux_output[2]~4_combout  = (always07 & (temp_aluResult_2)) # (!always07 & ((temp_rdat_one_output_2)))

	.dataa(temp_aluResult_2),
	.datab(gnd),
	.datac(temp_rdat_one_output_2),
	.datad(always03),
	.cin(gnd),
	.combout(\alu_a_mux_output[2]~4_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[2]~4 .lut_mask = 16'hAAF0;
defparam \alu_a_mux_output[2]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N10
cycloneive_lcell_comb \alu_a_mux_output[4]~6 (
// Equation(s):
// \alu_a_mux_output[4]~6_combout  = (always07 & ((temp_aluResult_4))) # (!always07 & (temp_rdat_one_output_4))

	.dataa(gnd),
	.datab(temp_rdat_one_output_4),
	.datac(temp_aluResult_4),
	.datad(always03),
	.cin(gnd),
	.combout(\alu_a_mux_output[4]~6_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[4]~6 .lut_mask = 16'hF0CC;
defparam \alu_a_mux_output[4]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N18
cycloneive_lcell_comb \alu_a_mux_output[8]~10 (
// Equation(s):
// \alu_a_mux_output[8]~10_combout  = (always07 & (temp_aluResult_8 & ((!forwarda_1)))) # (!always07 & (((Mux23 & forwarda_1))))

	.dataa(temp_aluResult_8),
	.datab(always03),
	.datac(Mux23),
	.datad(forwarda_1),
	.cin(gnd),
	.combout(\alu_a_mux_output[8]~10_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[8]~10 .lut_mask = 16'h3088;
defparam \alu_a_mux_output[8]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N6
cycloneive_lcell_comb \alu_a_mux_output[7]~12 (
// Equation(s):
// \alu_a_mux_output[7]~12_combout  = (forwarda_1 & (((!always07 & Mux24)))) # (!forwarda_1 & (temp_aluResult_7 & (always07)))

	.dataa(forwarda_1),
	.datab(temp_aluResult_7),
	.datac(always03),
	.datad(Mux24),
	.cin(gnd),
	.combout(\alu_a_mux_output[7]~12_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[7]~12 .lut_mask = 16'h4A40;
defparam \alu_a_mux_output[7]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N0
cycloneive_lcell_comb \alu_a_mux_output[6]~14 (
// Equation(s):
// \alu_a_mux_output[6]~14_combout  = (forwarda_1 & (Mux25 & (!always07))) # (!forwarda_1 & (((always07 & temp_aluResult_6))))

	.dataa(forwarda_1),
	.datab(Mux25),
	.datac(always03),
	.datad(temp_aluResult_6),
	.cin(gnd),
	.combout(\alu_a_mux_output[6]~14_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[6]~14 .lut_mask = 16'h5808;
defparam \alu_a_mux_output[6]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N12
cycloneive_lcell_comb \alu_a_mux_output[5]~16 (
// Equation(s):
// \alu_a_mux_output[5]~16_combout  = (always07 & (((temp_aluResult_5 & !forwarda_1)))) # (!always07 & (Mux26 & ((forwarda_1))))

	.dataa(always03),
	.datab(Mux26),
	.datac(temp_aluResult_5),
	.datad(forwarda_1),
	.cin(gnd),
	.combout(\alu_a_mux_output[5]~16_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[5]~16 .lut_mask = 16'h44A0;
defparam \alu_a_mux_output[5]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N14
cycloneive_lcell_comb \alu_a_mux_output[16]~18 (
// Equation(s):
// \alu_a_mux_output[16]~18_combout  = (always04) # ((!always07 & ((!always01) # (!always05))))

	.dataa(always02),
	.datab(always0),
	.datac(always03),
	.datad(always01),
	.cin(gnd),
	.combout(\alu_a_mux_output[16]~18_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[16]~18 .lut_mask = 16'hFF07;
defparam \alu_a_mux_output[16]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N0
cycloneive_lcell_comb \alu_a_mux_output[16]~19 (
// Equation(s):
// \alu_a_mux_output[16]~19_combout  = (forwarda_1 & ((\alu_a_mux_output[16]~18_combout ) # ((Mux15)))) # (!forwarda_1 & (!\alu_a_mux_output[16]~18_combout  & ((temp_aluResult_16))))

	.dataa(forwarda_1),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(Mux15),
	.datad(temp_aluResult_16),
	.cin(gnd),
	.combout(\alu_a_mux_output[16]~19_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[16]~19 .lut_mask = 16'hB9A8;
defparam \alu_a_mux_output[16]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N22
cycloneive_lcell_comb \alu_a_mux_output[14]~21 (
// Equation(s):
// \alu_a_mux_output[14]~21_combout  = (always07 & (temp_aluResult_14 & (!forwarda_1))) # (!always07 & (((forwarda_1 & Mux17))))

	.dataa(temp_aluResult_14),
	.datab(always03),
	.datac(forwarda_1),
	.datad(Mux17),
	.cin(gnd),
	.combout(\alu_a_mux_output[14]~21_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[14]~21 .lut_mask = 16'h3808;
defparam \alu_a_mux_output[14]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N12
cycloneive_lcell_comb \alu_a_mux_output[15]~23 (
// Equation(s):
// \alu_a_mux_output[15]~23_combout  = (forwarda_1 & (Mux16 & (!always07))) # (!forwarda_1 & (((always07 & temp_aluResult_15))))

	.dataa(Mux16),
	.datab(forwarda_1),
	.datac(always03),
	.datad(temp_aluResult_15),
	.cin(gnd),
	.combout(\alu_a_mux_output[15]~23_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[15]~23 .lut_mask = 16'h3808;
defparam \alu_a_mux_output[15]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N4
cycloneive_lcell_comb \alu_a_mux_output[13]~25 (
// Equation(s):
// \alu_a_mux_output[13]~25_combout  = (always07 & (temp_aluResult_13 & ((!forwarda_1)))) # (!always07 & (((Mux18 & forwarda_1))))

	.dataa(temp_aluResult_13),
	.datab(Mux18),
	.datac(always03),
	.datad(forwarda_1),
	.cin(gnd),
	.combout(\alu_a_mux_output[13]~25_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[13]~25 .lut_mask = 16'h0CA0;
defparam \alu_a_mux_output[13]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N30
cycloneive_lcell_comb \alu_a_mux_output[12]~27 (
// Equation(s):
// \alu_a_mux_output[12]~27_combout  = (forwarda_1 & (Mux19 & ((!always07)))) # (!forwarda_1 & (((temp_aluResult_12 & always07))))

	.dataa(Mux19),
	.datab(forwarda_1),
	.datac(temp_aluResult_12),
	.datad(always03),
	.cin(gnd),
	.combout(\alu_a_mux_output[12]~27_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[12]~27 .lut_mask = 16'h3088;
defparam \alu_a_mux_output[12]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N12
cycloneive_lcell_comb \alu_a_mux_output[10]~29 (
// Equation(s):
// \alu_a_mux_output[10]~29_combout  = (forwarda_1 & (!always07 & ((Mux21)))) # (!forwarda_1 & (always07 & (temp_aluResult_10)))

	.dataa(forwarda_1),
	.datab(always03),
	.datac(temp_aluResult_10),
	.datad(Mux21),
	.cin(gnd),
	.combout(\alu_a_mux_output[10]~29_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[10]~29 .lut_mask = 16'h6240;
defparam \alu_a_mux_output[10]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N0
cycloneive_lcell_comb \alu_a_mux_output[11]~31 (
// Equation(s):
// \alu_a_mux_output[11]~31_combout  = (always07 & (temp_aluResult_11 & ((!forwarda_1)))) # (!always07 & (((Mux20 & forwarda_1))))

	.dataa(temp_aluResult_11),
	.datab(always03),
	.datac(Mux20),
	.datad(forwarda_1),
	.cin(gnd),
	.combout(\alu_a_mux_output[11]~31_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[11]~31 .lut_mask = 16'h3088;
defparam \alu_a_mux_output[11]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N8
cycloneive_lcell_comb \alu_a_mux_output[9]~33 (
// Equation(s):
// \alu_a_mux_output[9]~33_combout  = (always07 & (((temp_aluResult_9 & !forwarda_1)))) # (!always07 & (Mux22 & ((forwarda_1))))

	.dataa(Mux22),
	.datab(temp_aluResult_9),
	.datac(always03),
	.datad(forwarda_1),
	.cin(gnd),
	.combout(\alu_a_mux_output[9]~33_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[9]~33 .lut_mask = 16'h0AC0;
defparam \alu_a_mux_output[9]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N22
cycloneive_lcell_comb \alu_a_mux_output[31]~35 (
// Equation(s):
// \alu_a_mux_output[31]~35_combout  = (\alu_a_mux_output[16]~18_combout  & (forwarda_1)) # (!\alu_a_mux_output[16]~18_combout  & ((forwarda_1 & ((Mux0))) # (!forwarda_1 & (temp_aluResult_31))))

	.dataa(\alu_a_mux_output[16]~18_combout ),
	.datab(forwarda_1),
	.datac(temp_aluResult_31),
	.datad(Mux0),
	.cin(gnd),
	.combout(\alu_a_mux_output[31]~35_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[31]~35 .lut_mask = 16'hDC98;
defparam \alu_a_mux_output[31]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N28
cycloneive_lcell_comb \alu_a_mux_output[30]~37 (
// Equation(s):
// \alu_a_mux_output[30]~37_combout  = (\alu_a_mux_output[16]~18_combout  & (forwarda_1)) # (!\alu_a_mux_output[16]~18_combout  & ((forwarda_1 & (Mux1)) # (!forwarda_1 & ((temp_aluResult_30)))))

	.dataa(\alu_a_mux_output[16]~18_combout ),
	.datab(forwarda_1),
	.datac(Mux1),
	.datad(temp_aluResult_30),
	.cin(gnd),
	.combout(\alu_a_mux_output[30]~37_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[30]~37 .lut_mask = 16'hD9C8;
defparam \alu_a_mux_output[30]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N26
cycloneive_lcell_comb \alu_a_mux_output[29]~39 (
// Equation(s):
// \alu_a_mux_output[29]~39_combout  = (forwarda_1 & ((Mux2) # ((\alu_a_mux_output[16]~18_combout )))) # (!forwarda_1 & (((!\alu_a_mux_output[16]~18_combout  & temp_aluResult_29))))

	.dataa(Mux2),
	.datab(forwarda_1),
	.datac(\alu_a_mux_output[16]~18_combout ),
	.datad(temp_aluResult_29),
	.cin(gnd),
	.combout(\alu_a_mux_output[29]~39_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[29]~39 .lut_mask = 16'hCBC8;
defparam \alu_a_mux_output[29]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N18
cycloneive_lcell_comb \alu_a_mux_output[26]~41 (
// Equation(s):
// \alu_a_mux_output[26]~41_combout  = (\alu_a_mux_output[16]~18_combout  & (((forwarda_1)))) # (!\alu_a_mux_output[16]~18_combout  & ((forwarda_1 & (Mux5)) # (!forwarda_1 & ((temp_aluResult_26)))))

	.dataa(Mux5),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(temp_aluResult_26),
	.datad(forwarda_1),
	.cin(gnd),
	.combout(\alu_a_mux_output[26]~41_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[26]~41 .lut_mask = 16'hEE30;
defparam \alu_a_mux_output[26]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N12
cycloneive_lcell_comb \alu_a_mux_output[25]~43 (
// Equation(s):
// \alu_a_mux_output[25]~43_combout  = (forwarda_1 & (((\alu_a_mux_output[16]~18_combout ) # (Mux6)))) # (!forwarda_1 & (temp_aluResult_25 & (!\alu_a_mux_output[16]~18_combout )))

	.dataa(forwarda_1),
	.datab(temp_aluResult_25),
	.datac(\alu_a_mux_output[16]~18_combout ),
	.datad(Mux6),
	.cin(gnd),
	.combout(\alu_a_mux_output[25]~43_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[25]~43 .lut_mask = 16'hAEA4;
defparam \alu_a_mux_output[25]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N14
cycloneive_lcell_comb \alu_a_mux_output[28]~45 (
// Equation(s):
// \alu_a_mux_output[28]~45_combout  = (\alu_a_mux_output[16]~18_combout  & (((forwarda_1)))) # (!\alu_a_mux_output[16]~18_combout  & ((forwarda_1 & (Mux3)) # (!forwarda_1 & ((temp_aluResult_28)))))

	.dataa(Mux3),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(forwarda_1),
	.datad(temp_aluResult_28),
	.cin(gnd),
	.combout(\alu_a_mux_output[28]~45_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[28]~45 .lut_mask = 16'hE3E0;
defparam \alu_a_mux_output[28]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N22
cycloneive_lcell_comb \alu_a_mux_output[27]~47 (
// Equation(s):
// \alu_a_mux_output[27]~47_combout  = (\alu_a_mux_output[16]~18_combout  & (forwarda_1)) # (!\alu_a_mux_output[16]~18_combout  & ((forwarda_1 & (Mux4)) # (!forwarda_1 & ((temp_aluResult_27)))))

	.dataa(\alu_a_mux_output[16]~18_combout ),
	.datab(forwarda_1),
	.datac(Mux4),
	.datad(temp_aluResult_27),
	.cin(gnd),
	.combout(\alu_a_mux_output[27]~47_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[27]~47 .lut_mask = 16'hD9C8;
defparam \alu_a_mux_output[27]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N30
cycloneive_lcell_comb \alu_a_mux_output[17]~49 (
// Equation(s):
// \alu_a_mux_output[17]~49_combout  = (forwarda_1 & ((Mux14) # ((\alu_a_mux_output[16]~18_combout )))) # (!forwarda_1 & (((temp_aluResult_17 & !\alu_a_mux_output[16]~18_combout ))))

	.dataa(forwarda_1),
	.datab(Mux14),
	.datac(temp_aluResult_17),
	.datad(\alu_a_mux_output[16]~18_combout ),
	.cin(gnd),
	.combout(\alu_a_mux_output[17]~49_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[17]~49 .lut_mask = 16'hAAD8;
defparam \alu_a_mux_output[17]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N18
cycloneive_lcell_comb \alu_a_mux_output[20]~51 (
// Equation(s):
// \alu_a_mux_output[20]~51_combout  = (forwarda_1 & ((Mux11) # ((\alu_a_mux_output[16]~18_combout )))) # (!forwarda_1 & (((temp_aluResult_20 & !\alu_a_mux_output[16]~18_combout ))))

	.dataa(Mux11),
	.datab(temp_aluResult_20),
	.datac(forwarda_1),
	.datad(\alu_a_mux_output[16]~18_combout ),
	.cin(gnd),
	.combout(\alu_a_mux_output[20]~51_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[20]~51 .lut_mask = 16'hF0AC;
defparam \alu_a_mux_output[20]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N20
cycloneive_lcell_comb \alu_a_mux_output[19]~53 (
// Equation(s):
// \alu_a_mux_output[19]~53_combout  = (\alu_a_mux_output[16]~18_combout  & (((forwarda_1)))) # (!\alu_a_mux_output[16]~18_combout  & ((forwarda_1 & (Mux12)) # (!forwarda_1 & ((temp_aluResult_19)))))

	.dataa(Mux12),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(forwarda_1),
	.datad(temp_aluResult_19),
	.cin(gnd),
	.combout(\alu_a_mux_output[19]~53_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[19]~53 .lut_mask = 16'hE3E0;
defparam \alu_a_mux_output[19]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N20
cycloneive_lcell_comb \alu_a_mux_output[18]~55 (
// Equation(s):
// \alu_a_mux_output[18]~55_combout  = (\alu_a_mux_output[16]~18_combout  & (forwarda_1)) # (!\alu_a_mux_output[16]~18_combout  & ((forwarda_1 & (Mux13)) # (!forwarda_1 & ((temp_aluResult_18)))))

	.dataa(\alu_a_mux_output[16]~18_combout ),
	.datab(forwarda_1),
	.datac(Mux13),
	.datad(temp_aluResult_18),
	.cin(gnd),
	.combout(\alu_a_mux_output[18]~55_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[18]~55 .lut_mask = 16'hD9C8;
defparam \alu_a_mux_output[18]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N6
cycloneive_lcell_comb \alu_a_mux_output[24]~57 (
// Equation(s):
// \alu_a_mux_output[24]~57_combout  = (forwarda_1 & ((\alu_a_mux_output[16]~18_combout ) # ((Mux7)))) # (!forwarda_1 & (!\alu_a_mux_output[16]~18_combout  & (temp_aluResult_24)))

	.dataa(forwarda_1),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(temp_aluResult_24),
	.datad(Mux7),
	.cin(gnd),
	.combout(\alu_a_mux_output[24]~57_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[24]~57 .lut_mask = 16'hBA98;
defparam \alu_a_mux_output[24]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N16
cycloneive_lcell_comb \alu_a_mux_output[23]~59 (
// Equation(s):
// \alu_a_mux_output[23]~59_combout  = (forwarda_1 & ((\alu_a_mux_output[16]~18_combout ) # ((Mux8)))) # (!forwarda_1 & (!\alu_a_mux_output[16]~18_combout  & (temp_aluResult_23)))

	.dataa(forwarda_1),
	.datab(\alu_a_mux_output[16]~18_combout ),
	.datac(temp_aluResult_23),
	.datad(Mux8),
	.cin(gnd),
	.combout(\alu_a_mux_output[23]~59_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[23]~59 .lut_mask = 16'hBA98;
defparam \alu_a_mux_output[23]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N16
cycloneive_lcell_comb \alu_a_mux_output[22]~61 (
// Equation(s):
// \alu_a_mux_output[22]~61_combout  = (forwarda_1 & ((Mux9) # ((\alu_a_mux_output[16]~18_combout )))) # (!forwarda_1 & (((temp_aluResult_22 & !\alu_a_mux_output[16]~18_combout ))))

	.dataa(Mux9),
	.datab(temp_aluResult_22),
	.datac(forwarda_1),
	.datad(\alu_a_mux_output[16]~18_combout ),
	.cin(gnd),
	.combout(\alu_a_mux_output[22]~61_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[22]~61 .lut_mask = 16'hF0AC;
defparam \alu_a_mux_output[22]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N20
cycloneive_lcell_comb \alu_a_mux_output[21]~63 (
// Equation(s):
// \alu_a_mux_output[21]~63_combout  = (forwarda_1 & (((Mux10) # (\alu_a_mux_output[16]~18_combout )))) # (!forwarda_1 & (temp_aluResult_21 & ((!\alu_a_mux_output[16]~18_combout ))))

	.dataa(forwarda_1),
	.datab(temp_aluResult_21),
	.datac(Mux10),
	.datad(\alu_a_mux_output[16]~18_combout ),
	.cin(gnd),
	.combout(\alu_a_mux_output[21]~63_combout ),
	.cout());
// synopsys translate_off
defparam \alu_a_mux_output[21]~63 .lut_mask = 16'hAAE4;
defparam \alu_a_mux_output[21]~63 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module alu_b_mux (
	temp_aluResult_1,
	temp_aluResult_0,
	temp_aluResult_2,
	temp_aluResult_3,
	temp_aluResult_5,
	temp_aluResult_4,
	temp_aluResult_7,
	temp_aluResult_6,
	temp_aluResult_9,
	temp_aluResult_8,
	temp_aluResult_11,
	temp_aluResult_10,
	temp_aluResult_13,
	temp_aluResult_12,
	temp_aluResult_15,
	temp_aluResult_14,
	temp_aluResult_17,
	temp_aluResult_16,
	temp_aluResult_19,
	temp_aluResult_18,
	temp_aluResult_20,
	temp_aluResult_21,
	temp_aluResult_23,
	temp_aluResult_22,
	temp_aluResult_25,
	temp_aluResult_24,
	temp_aluResult_26,
	temp_aluResult_27,
	temp_aluResult_29,
	temp_aluResult_28,
	temp_aluResult_31,
	temp_aluResult_30,
	temp_rdat_two_output_1,
	always0,
	always01,
	always02,
	alu_b_mux_output_1,
	Mux30,
	always03,
	forwardb_1,
	alu_b_mux_output_11,
	Mux31,
	alu_b_mux_output_0,
	temp_rdat_two_output_0,
	alu_b_mux_output_01,
	Mux29,
	Mux27,
	Mux28,
	temp_rdat_two_output_2,
	alu_b_mux_output_2,
	Mux23,
	Mux24,
	Mux25,
	Mux26,
	temp_rdat_two_output_3,
	alu_b_mux_output_3,
	Mux15,
	temp_iMemLoad_0,
	Mux17,
	Mux16,
	Mux18,
	Mux19,
	Mux21,
	Mux20,
	Mux22,
	temp_rdat_two_output_4,
	alu_b_mux_output_4,
	Mux0,
	temp_iMemLoad_15,
	Mux1,
	temp_iMemLoad_14,
	Mux2,
	temp_iMemLoad_13,
	Mux5,
	temp_iMemLoad_10,
	Mux6,
	temp_iMemLoad_9,
	Mux3,
	temp_iMemLoad_12,
	Mux4,
	temp_iMemLoad_11,
	Mux14,
	temp_iMemLoad_1,
	Mux11,
	temp_iMemLoad_4,
	Mux12,
	temp_iMemLoad_3,
	Mux13,
	temp_iMemLoad_2,
	Mux7,
	temp_iMemLoad_8,
	Mux8,
	temp_iMemLoad_7,
	Mux9,
	temp_iMemLoad_6,
	Mux10,
	temp_iMemLoad_5,
	temp_rdat_two_output_15,
	alu_b_mux_output_15,
	temp_rdat_two_output_12,
	alu_b_mux_output_12,
	temp_rdat_two_output_27,
	alu_b_mux_output_27,
	temp_rdat_two_output_18,
	alu_b_mux_output_18,
	temp_rdat_two_output_17,
	alu_b_mux_output_17,
	temp_rdat_two_output_16,
	alu_b_mux_output_16,
	temp_rdat_two_output_31,
	alu_b_mux_output_31,
	temp_rdat_two_output_30,
	alu_b_mux_output_30,
	temp_rdat_two_output_29,
	alu_b_mux_output_29,
	temp_rdat_two_output_28,
	alu_b_mux_output_28,
	temp_rdat_two_output_26,
	alu_b_mux_output_26,
	temp_rdat_two_output_25,
	alu_b_mux_output_25,
	temp_rdat_two_output_24,
	alu_b_mux_output_24,
	temp_rdat_two_output_23,
	alu_b_mux_output_23,
	temp_rdat_two_output_22,
	alu_b_mux_output_22,
	temp_rdat_two_output_21,
	alu_b_mux_output_21,
	temp_rdat_two_output_20,
	alu_b_mux_output_20,
	temp_rdat_two_output_19,
	alu_b_mux_output_19,
	temp_rdat_two_output_10,
	alu_b_mux_output_10,
	temp_rdat_two_output_14,
	alu_b_mux_output_14,
	temp_rdat_two_output_9,
	alu_b_mux_output_9,
	temp_rdat_two_output_8,
	alu_b_mux_output_8,
	temp_rdat_two_output_7,
	alu_b_mux_output_7,
	temp_rdat_two_output_6,
	alu_b_mux_output_6,
	temp_rdat_two_output_5,
	alu_b_mux_output_5,
	temp_rdat_two_output_13,
	alu_b_mux_output_13,
	temp_rdat_two_output_11,
	alu_b_mux_output_111,
	always04,
	devpor,
	devclrn,
	devoe);
input 	temp_aluResult_1;
input 	temp_aluResult_0;
input 	temp_aluResult_2;
input 	temp_aluResult_3;
input 	temp_aluResult_5;
input 	temp_aluResult_4;
input 	temp_aluResult_7;
input 	temp_aluResult_6;
input 	temp_aluResult_9;
input 	temp_aluResult_8;
input 	temp_aluResult_11;
input 	temp_aluResult_10;
input 	temp_aluResult_13;
input 	temp_aluResult_12;
input 	temp_aluResult_15;
input 	temp_aluResult_14;
input 	temp_aluResult_17;
input 	temp_aluResult_16;
input 	temp_aluResult_19;
input 	temp_aluResult_18;
input 	temp_aluResult_20;
input 	temp_aluResult_21;
input 	temp_aluResult_23;
input 	temp_aluResult_22;
input 	temp_aluResult_25;
input 	temp_aluResult_24;
input 	temp_aluResult_26;
input 	temp_aluResult_27;
input 	temp_aluResult_29;
input 	temp_aluResult_28;
input 	temp_aluResult_31;
input 	temp_aluResult_30;
input 	temp_rdat_two_output_1;
input 	always0;
input 	always01;
input 	always02;
output 	alu_b_mux_output_1;
input 	Mux30;
input 	always03;
input 	forwardb_1;
output 	alu_b_mux_output_11;
input 	Mux31;
output 	alu_b_mux_output_0;
input 	temp_rdat_two_output_0;
output 	alu_b_mux_output_01;
input 	Mux29;
input 	Mux27;
input 	Mux28;
input 	temp_rdat_two_output_2;
output 	alu_b_mux_output_2;
input 	Mux23;
input 	Mux24;
input 	Mux25;
input 	Mux26;
input 	temp_rdat_two_output_3;
output 	alu_b_mux_output_3;
input 	Mux15;
input 	temp_iMemLoad_0;
input 	Mux17;
input 	Mux16;
input 	Mux18;
input 	Mux19;
input 	Mux21;
input 	Mux20;
input 	Mux22;
input 	temp_rdat_two_output_4;
output 	alu_b_mux_output_4;
input 	Mux0;
input 	temp_iMemLoad_15;
input 	Mux1;
input 	temp_iMemLoad_14;
input 	Mux2;
input 	temp_iMemLoad_13;
input 	Mux5;
input 	temp_iMemLoad_10;
input 	Mux6;
input 	temp_iMemLoad_9;
input 	Mux3;
input 	temp_iMemLoad_12;
input 	Mux4;
input 	temp_iMemLoad_11;
input 	Mux14;
input 	temp_iMemLoad_1;
input 	Mux11;
input 	temp_iMemLoad_4;
input 	Mux12;
input 	temp_iMemLoad_3;
input 	Mux13;
input 	temp_iMemLoad_2;
input 	Mux7;
input 	temp_iMemLoad_8;
input 	Mux8;
input 	temp_iMemLoad_7;
input 	Mux9;
input 	temp_iMemLoad_6;
input 	Mux10;
input 	temp_iMemLoad_5;
input 	temp_rdat_two_output_15;
output 	alu_b_mux_output_15;
input 	temp_rdat_two_output_12;
output 	alu_b_mux_output_12;
input 	temp_rdat_two_output_27;
output 	alu_b_mux_output_27;
input 	temp_rdat_two_output_18;
output 	alu_b_mux_output_18;
input 	temp_rdat_two_output_17;
output 	alu_b_mux_output_17;
input 	temp_rdat_two_output_16;
output 	alu_b_mux_output_16;
input 	temp_rdat_two_output_31;
output 	alu_b_mux_output_31;
input 	temp_rdat_two_output_30;
output 	alu_b_mux_output_30;
input 	temp_rdat_two_output_29;
output 	alu_b_mux_output_29;
input 	temp_rdat_two_output_28;
output 	alu_b_mux_output_28;
input 	temp_rdat_two_output_26;
output 	alu_b_mux_output_26;
input 	temp_rdat_two_output_25;
output 	alu_b_mux_output_25;
input 	temp_rdat_two_output_24;
output 	alu_b_mux_output_24;
input 	temp_rdat_two_output_23;
output 	alu_b_mux_output_23;
input 	temp_rdat_two_output_22;
output 	alu_b_mux_output_22;
input 	temp_rdat_two_output_21;
output 	alu_b_mux_output_21;
input 	temp_rdat_two_output_20;
output 	alu_b_mux_output_20;
input 	temp_rdat_two_output_19;
output 	alu_b_mux_output_19;
input 	temp_rdat_two_output_10;
output 	alu_b_mux_output_10;
input 	temp_rdat_two_output_14;
output 	alu_b_mux_output_14;
input 	temp_rdat_two_output_9;
output 	alu_b_mux_output_9;
input 	temp_rdat_two_output_8;
output 	alu_b_mux_output_8;
input 	temp_rdat_two_output_7;
output 	alu_b_mux_output_7;
input 	temp_rdat_two_output_6;
output 	alu_b_mux_output_6;
input 	temp_rdat_two_output_5;
output 	alu_b_mux_output_5;
input 	temp_rdat_two_output_13;
output 	alu_b_mux_output_13;
input 	temp_rdat_two_output_11;
output 	alu_b_mux_output_111;
input 	always04;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \alu_b_mux_output[2]~4_combout ;
wire \alu_b_mux_output[3]~6_combout ;
wire \alu_b_mux_output[4]~8_combout ;
wire \alu_b_mux_output[15]~10_combout ;
wire \alu_b_mux_output[12]~12_combout ;
wire \alu_b_mux_output[27]~14_combout ;
wire \alu_b_mux_output[27]~15_combout ;
wire \alu_b_mux_output[18]~17_combout ;
wire \alu_b_mux_output[17]~19_combout ;
wire \alu_b_mux_output[16]~21_combout ;
wire \alu_b_mux_output[31]~23_combout ;
wire \alu_b_mux_output[30]~25_combout ;
wire \alu_b_mux_output[29]~27_combout ;
wire \alu_b_mux_output[28]~29_combout ;
wire \alu_b_mux_output[26]~31_combout ;
wire \alu_b_mux_output[25]~33_combout ;
wire \alu_b_mux_output[24]~35_combout ;
wire \alu_b_mux_output[23]~37_combout ;
wire \alu_b_mux_output[22]~39_combout ;
wire \alu_b_mux_output[21]~41_combout ;
wire \alu_b_mux_output[20]~43_combout ;
wire \alu_b_mux_output[19]~45_combout ;
wire \alu_b_mux_output[10]~47_combout ;
wire \alu_b_mux_output[14]~49_combout ;
wire \alu_b_mux_output[9]~51_combout ;
wire \alu_b_mux_output[8]~53_combout ;
wire \alu_b_mux_output[7]~55_combout ;
wire \alu_b_mux_output[6]~57_combout ;
wire \alu_b_mux_output[5]~59_combout ;
wire \alu_b_mux_output[13]~61_combout ;
wire \alu_b_mux_output[11]~63_combout ;


// Location: LCCOMB_X61_Y39_N20
cycloneive_lcell_comb \alu_b_mux_output[1]~0 (
// Equation(s):
// alu_b_mux_output_1 = (!always06 & (temp_rdat_two_output_1 & (!always02 & !always0)))

	.dataa(always04),
	.datab(temp_rdat_two_output_1),
	.datac(always02),
	.datad(always0),
	.cin(gnd),
	.combout(alu_b_mux_output_1),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[1]~0 .lut_mask = 16'h0004;
defparam \alu_b_mux_output[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N16
cycloneive_lcell_comb \alu_b_mux_output[1]~1 (
// Equation(s):
// alu_b_mux_output_11 = (always06 & (temp_aluResult_1 & (!forwardb_1))) # (!always06 & (((forwardb_1 & Mux30))))

	.dataa(temp_aluResult_1),
	.datab(always04),
	.datac(forwardb_1),
	.datad(Mux30),
	.cin(gnd),
	.combout(alu_b_mux_output_11),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[1]~1 .lut_mask = 16'h3808;
defparam \alu_b_mux_output[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N30
cycloneive_lcell_comb \alu_b_mux_output[0]~2 (
// Equation(s):
// alu_b_mux_output_0 = (forwardb_1 & (Mux31 & (!always06))) # (!forwardb_1 & (((always06 & temp_aluResult_0))))

	.dataa(forwardb_1),
	.datab(Mux31),
	.datac(always04),
	.datad(temp_aluResult_0),
	.cin(gnd),
	.combout(alu_b_mux_output_0),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[0]~2 .lut_mask = 16'h5808;
defparam \alu_b_mux_output[0]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N2
cycloneive_lcell_comb \alu_b_mux_output[0]~3 (
// Equation(s):
// alu_b_mux_output_01 = (!always06 & (temp_rdat_two_output_0 & (!always02 & !always0)))

	.dataa(always04),
	.datab(temp_rdat_two_output_0),
	.datac(always02),
	.datad(always0),
	.cin(gnd),
	.combout(alu_b_mux_output_01),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[0]~3 .lut_mask = 16'h0004;
defparam \alu_b_mux_output[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N18
cycloneive_lcell_comb \alu_b_mux_output[2]~5 (
// Equation(s):
// alu_b_mux_output_2 = (\alu_b_mux_output[2]~4_combout ) # ((!forwardb_1 & (temp_rdat_two_output_2 & !always06)))

	.dataa(forwardb_1),
	.datab(temp_rdat_two_output_2),
	.datac(always04),
	.datad(\alu_b_mux_output[2]~4_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_2),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[2]~5 .lut_mask = 16'hFF04;
defparam \alu_b_mux_output[2]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N14
cycloneive_lcell_comb \alu_b_mux_output[3]~7 (
// Equation(s):
// alu_b_mux_output_3 = (\alu_b_mux_output[3]~6_combout ) # ((!forwardb_1 & (temp_rdat_two_output_3 & !always06)))

	.dataa(forwardb_1),
	.datab(temp_rdat_two_output_3),
	.datac(\alu_b_mux_output[3]~6_combout ),
	.datad(always04),
	.cin(gnd),
	.combout(alu_b_mux_output_3),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[3]~7 .lut_mask = 16'hF0F4;
defparam \alu_b_mux_output[3]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N28
cycloneive_lcell_comb \alu_b_mux_output[4]~9 (
// Equation(s):
// alu_b_mux_output_4 = (\alu_b_mux_output[4]~8_combout ) # ((temp_rdat_two_output_4 & (!forwardb_1 & !always06)))

	.dataa(temp_rdat_two_output_4),
	.datab(\alu_b_mux_output[4]~8_combout ),
	.datac(forwardb_1),
	.datad(always04),
	.cin(gnd),
	.combout(alu_b_mux_output_4),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[4]~9 .lut_mask = 16'hCCCE;
defparam \alu_b_mux_output[4]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N8
cycloneive_lcell_comb \alu_b_mux_output[15]~11 (
// Equation(s):
// alu_b_mux_output_15 = (\alu_b_mux_output[15]~10_combout ) # ((!forwardb_1 & (temp_rdat_two_output_15 & !always06)))

	.dataa(forwardb_1),
	.datab(temp_rdat_two_output_15),
	.datac(\alu_b_mux_output[15]~10_combout ),
	.datad(always04),
	.cin(gnd),
	.combout(alu_b_mux_output_15),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[15]~11 .lut_mask = 16'hF0F4;
defparam \alu_b_mux_output[15]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N2
cycloneive_lcell_comb \alu_b_mux_output[12]~13 (
// Equation(s):
// alu_b_mux_output_12 = (\alu_b_mux_output[12]~12_combout ) # ((!always06 & (temp_rdat_two_output_12 & !forwardb_1)))

	.dataa(\alu_b_mux_output[12]~12_combout ),
	.datab(always04),
	.datac(temp_rdat_two_output_12),
	.datad(forwardb_1),
	.cin(gnd),
	.combout(alu_b_mux_output_12),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[12]~13 .lut_mask = 16'hAABA;
defparam \alu_b_mux_output[12]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N24
cycloneive_lcell_comb \alu_b_mux_output[27]~16 (
// Equation(s):
// alu_b_mux_output_27 = (\alu_b_mux_output[27]~14_combout  & ((\alu_b_mux_output[27]~15_combout  & ((temp_iMemLoad_11))) # (!\alu_b_mux_output[27]~15_combout  & (temp_rdat_two_output_27)))) # (!\alu_b_mux_output[27]~14_combout  & 
// (((\alu_b_mux_output[27]~15_combout ))))

	.dataa(temp_rdat_two_output_27),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(temp_iMemLoad_11),
	.datad(\alu_b_mux_output[27]~15_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_27),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[27]~16 .lut_mask = 16'hF388;
defparam \alu_b_mux_output[27]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N16
cycloneive_lcell_comb \alu_b_mux_output[18]~18 (
// Equation(s):
// alu_b_mux_output_18 = (\alu_b_mux_output[27]~14_combout  & ((\alu_b_mux_output[18]~17_combout  & (temp_iMemLoad_2)) # (!\alu_b_mux_output[18]~17_combout  & ((temp_rdat_two_output_18))))) # (!\alu_b_mux_output[27]~14_combout  & 
// (((\alu_b_mux_output[18]~17_combout ))))

	.dataa(temp_iMemLoad_2),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(temp_rdat_two_output_18),
	.datad(\alu_b_mux_output[18]~17_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_18),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[18]~18 .lut_mask = 16'hBBC0;
defparam \alu_b_mux_output[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N26
cycloneive_lcell_comb \alu_b_mux_output[17]~20 (
// Equation(s):
// alu_b_mux_output_17 = (\alu_b_mux_output[17]~19_combout  & (((temp_iMemLoad_1) # (!\alu_b_mux_output[27]~14_combout )))) # (!\alu_b_mux_output[17]~19_combout  & (temp_rdat_two_output_17 & (\alu_b_mux_output[27]~14_combout )))

	.dataa(temp_rdat_two_output_17),
	.datab(\alu_b_mux_output[17]~19_combout ),
	.datac(\alu_b_mux_output[27]~14_combout ),
	.datad(temp_iMemLoad_1),
	.cin(gnd),
	.combout(alu_b_mux_output_17),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[17]~20 .lut_mask = 16'hEC2C;
defparam \alu_b_mux_output[17]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N10
cycloneive_lcell_comb \alu_b_mux_output[16]~22 (
// Equation(s):
// alu_b_mux_output_16 = (\alu_b_mux_output[16]~21_combout  & ((temp_iMemLoad_0) # ((!\alu_b_mux_output[27]~14_combout )))) # (!\alu_b_mux_output[16]~21_combout  & (((temp_rdat_two_output_16 & \alu_b_mux_output[27]~14_combout ))))

	.dataa(temp_iMemLoad_0),
	.datab(temp_rdat_two_output_16),
	.datac(\alu_b_mux_output[16]~21_combout ),
	.datad(\alu_b_mux_output[27]~14_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_16),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[16]~22 .lut_mask = 16'hACF0;
defparam \alu_b_mux_output[16]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N12
cycloneive_lcell_comb \alu_b_mux_output[31]~24 (
// Equation(s):
// alu_b_mux_output_31 = (\alu_b_mux_output[27]~14_combout  & ((\alu_b_mux_output[31]~23_combout  & ((temp_iMemLoad_15))) # (!\alu_b_mux_output[31]~23_combout  & (temp_rdat_two_output_31)))) # (!\alu_b_mux_output[27]~14_combout  & 
// (((\alu_b_mux_output[31]~23_combout ))))

	.dataa(temp_rdat_two_output_31),
	.datab(temp_iMemLoad_15),
	.datac(\alu_b_mux_output[27]~14_combout ),
	.datad(\alu_b_mux_output[31]~23_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_31),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[31]~24 .lut_mask = 16'hCFA0;
defparam \alu_b_mux_output[31]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N26
cycloneive_lcell_comb \alu_b_mux_output[30]~26 (
// Equation(s):
// alu_b_mux_output_30 = (\alu_b_mux_output[27]~14_combout  & ((\alu_b_mux_output[30]~25_combout  & (temp_iMemLoad_14)) # (!\alu_b_mux_output[30]~25_combout  & ((temp_rdat_two_output_30))))) # (!\alu_b_mux_output[27]~14_combout  & 
// (((\alu_b_mux_output[30]~25_combout ))))

	.dataa(temp_iMemLoad_14),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(temp_rdat_two_output_30),
	.datad(\alu_b_mux_output[30]~25_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_30),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[30]~26 .lut_mask = 16'hBBC0;
defparam \alu_b_mux_output[30]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N20
cycloneive_lcell_comb \alu_b_mux_output[29]~28 (
// Equation(s):
// alu_b_mux_output_29 = (\alu_b_mux_output[27]~14_combout  & ((\alu_b_mux_output[29]~27_combout  & (temp_iMemLoad_13)) # (!\alu_b_mux_output[29]~27_combout  & ((temp_rdat_two_output_29))))) # (!\alu_b_mux_output[27]~14_combout  & 
// (((\alu_b_mux_output[29]~27_combout ))))

	.dataa(\alu_b_mux_output[27]~14_combout ),
	.datab(temp_iMemLoad_13),
	.datac(\alu_b_mux_output[29]~27_combout ),
	.datad(temp_rdat_two_output_29),
	.cin(gnd),
	.combout(alu_b_mux_output_29),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[29]~28 .lut_mask = 16'hDAD0;
defparam \alu_b_mux_output[29]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N24
cycloneive_lcell_comb \alu_b_mux_output[28]~30 (
// Equation(s):
// alu_b_mux_output_28 = (\alu_b_mux_output[27]~14_combout  & ((\alu_b_mux_output[28]~29_combout  & (temp_iMemLoad_12)) # (!\alu_b_mux_output[28]~29_combout  & ((temp_rdat_two_output_28))))) # (!\alu_b_mux_output[27]~14_combout  & 
// (((\alu_b_mux_output[28]~29_combout ))))

	.dataa(temp_iMemLoad_12),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(temp_rdat_two_output_28),
	.datad(\alu_b_mux_output[28]~29_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_28),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[28]~30 .lut_mask = 16'hBBC0;
defparam \alu_b_mux_output[28]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N0
cycloneive_lcell_comb \alu_b_mux_output[26]~32 (
// Equation(s):
// alu_b_mux_output_26 = (\alu_b_mux_output[27]~14_combout  & ((\alu_b_mux_output[26]~31_combout  & (temp_iMemLoad_10)) # (!\alu_b_mux_output[26]~31_combout  & ((temp_rdat_two_output_26))))) # (!\alu_b_mux_output[27]~14_combout  & 
// (((\alu_b_mux_output[26]~31_combout ))))

	.dataa(temp_iMemLoad_10),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(\alu_b_mux_output[26]~31_combout ),
	.datad(temp_rdat_two_output_26),
	.cin(gnd),
	.combout(alu_b_mux_output_26),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[26]~32 .lut_mask = 16'hBCB0;
defparam \alu_b_mux_output[26]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N28
cycloneive_lcell_comb \alu_b_mux_output[25]~34 (
// Equation(s):
// alu_b_mux_output_25 = (\alu_b_mux_output[25]~33_combout  & (((temp_iMemLoad_9) # (!\alu_b_mux_output[27]~14_combout )))) # (!\alu_b_mux_output[25]~33_combout  & (temp_rdat_two_output_25 & ((\alu_b_mux_output[27]~14_combout ))))

	.dataa(temp_rdat_two_output_25),
	.datab(temp_iMemLoad_9),
	.datac(\alu_b_mux_output[25]~33_combout ),
	.datad(\alu_b_mux_output[27]~14_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_25),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[25]~34 .lut_mask = 16'hCAF0;
defparam \alu_b_mux_output[25]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N12
cycloneive_lcell_comb \alu_b_mux_output[24]~36 (
// Equation(s):
// alu_b_mux_output_24 = (\alu_b_mux_output[27]~14_combout  & ((\alu_b_mux_output[24]~35_combout  & ((temp_iMemLoad_8))) # (!\alu_b_mux_output[24]~35_combout  & (temp_rdat_two_output_24)))) # (!\alu_b_mux_output[27]~14_combout  & 
// (((\alu_b_mux_output[24]~35_combout ))))

	.dataa(temp_rdat_two_output_24),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(temp_iMemLoad_8),
	.datad(\alu_b_mux_output[24]~35_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_24),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[24]~36 .lut_mask = 16'hF388;
defparam \alu_b_mux_output[24]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N0
cycloneive_lcell_comb \alu_b_mux_output[23]~38 (
// Equation(s):
// alu_b_mux_output_23 = (\alu_b_mux_output[23]~37_combout  & ((temp_iMemLoad_7) # ((!\alu_b_mux_output[27]~14_combout )))) # (!\alu_b_mux_output[23]~37_combout  & (((temp_rdat_two_output_23 & \alu_b_mux_output[27]~14_combout ))))

	.dataa(\alu_b_mux_output[23]~37_combout ),
	.datab(temp_iMemLoad_7),
	.datac(temp_rdat_two_output_23),
	.datad(\alu_b_mux_output[27]~14_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_23),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[23]~38 .lut_mask = 16'hD8AA;
defparam \alu_b_mux_output[23]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N26
cycloneive_lcell_comb \alu_b_mux_output[22]~40 (
// Equation(s):
// alu_b_mux_output_22 = (\alu_b_mux_output[27]~14_combout  & ((\alu_b_mux_output[22]~39_combout  & (temp_iMemLoad_6)) # (!\alu_b_mux_output[22]~39_combout  & ((temp_rdat_two_output_22))))) # (!\alu_b_mux_output[27]~14_combout  & 
// (((\alu_b_mux_output[22]~39_combout ))))

	.dataa(temp_iMemLoad_6),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(\alu_b_mux_output[22]~39_combout ),
	.datad(temp_rdat_two_output_22),
	.cin(gnd),
	.combout(alu_b_mux_output_22),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[22]~40 .lut_mask = 16'hBCB0;
defparam \alu_b_mux_output[22]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N28
cycloneive_lcell_comb \alu_b_mux_output[21]~42 (
// Equation(s):
// alu_b_mux_output_21 = (\alu_b_mux_output[27]~14_combout  & ((\alu_b_mux_output[21]~41_combout  & ((temp_iMemLoad_5))) # (!\alu_b_mux_output[21]~41_combout  & (temp_rdat_two_output_21)))) # (!\alu_b_mux_output[27]~14_combout  & 
// (((\alu_b_mux_output[21]~41_combout ))))

	.dataa(\alu_b_mux_output[27]~14_combout ),
	.datab(temp_rdat_two_output_21),
	.datac(temp_iMemLoad_5),
	.datad(\alu_b_mux_output[21]~41_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_21),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[21]~42 .lut_mask = 16'hF588;
defparam \alu_b_mux_output[21]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N28
cycloneive_lcell_comb \alu_b_mux_output[20]~44 (
// Equation(s):
// alu_b_mux_output_20 = (\alu_b_mux_output[20]~43_combout  & (((temp_iMemLoad_4)) # (!\alu_b_mux_output[27]~14_combout ))) # (!\alu_b_mux_output[20]~43_combout  & (\alu_b_mux_output[27]~14_combout  & ((temp_rdat_two_output_20))))

	.dataa(\alu_b_mux_output[20]~43_combout ),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(temp_iMemLoad_4),
	.datad(temp_rdat_two_output_20),
	.cin(gnd),
	.combout(alu_b_mux_output_20),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[20]~44 .lut_mask = 16'hE6A2;
defparam \alu_b_mux_output[20]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N20
cycloneive_lcell_comb \alu_b_mux_output[19]~46 (
// Equation(s):
// alu_b_mux_output_19 = (\alu_b_mux_output[19]~45_combout  & (((temp_iMemLoad_3) # (!\alu_b_mux_output[27]~14_combout )))) # (!\alu_b_mux_output[19]~45_combout  & (temp_rdat_two_output_19 & ((\alu_b_mux_output[27]~14_combout ))))

	.dataa(\alu_b_mux_output[19]~45_combout ),
	.datab(temp_rdat_two_output_19),
	.datac(temp_iMemLoad_3),
	.datad(\alu_b_mux_output[27]~14_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_19),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[19]~46 .lut_mask = 16'hE4AA;
defparam \alu_b_mux_output[19]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N2
cycloneive_lcell_comb \alu_b_mux_output[10]~48 (
// Equation(s):
// alu_b_mux_output_10 = (\alu_b_mux_output[10]~47_combout ) # ((!forwardb_1 & (!always06 & temp_rdat_two_output_10)))

	.dataa(forwardb_1),
	.datab(always04),
	.datac(\alu_b_mux_output[10]~47_combout ),
	.datad(temp_rdat_two_output_10),
	.cin(gnd),
	.combout(alu_b_mux_output_10),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[10]~48 .lut_mask = 16'hF1F0;
defparam \alu_b_mux_output[10]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N14
cycloneive_lcell_comb \alu_b_mux_output[14]~50 (
// Equation(s):
// alu_b_mux_output_14 = (\alu_b_mux_output[14]~49_combout ) # ((temp_rdat_two_output_14 & (!always06 & !forwardb_1)))

	.dataa(temp_rdat_two_output_14),
	.datab(always04),
	.datac(forwardb_1),
	.datad(\alu_b_mux_output[14]~49_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_14),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[14]~50 .lut_mask = 16'hFF02;
defparam \alu_b_mux_output[14]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N14
cycloneive_lcell_comb \alu_b_mux_output[9]~52 (
// Equation(s):
// alu_b_mux_output_9 = (\alu_b_mux_output[9]~51_combout ) # ((!forwardb_1 & (!always06 & temp_rdat_two_output_9)))

	.dataa(forwardb_1),
	.datab(\alu_b_mux_output[9]~51_combout ),
	.datac(always04),
	.datad(temp_rdat_two_output_9),
	.cin(gnd),
	.combout(alu_b_mux_output_9),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[9]~52 .lut_mask = 16'hCDCC;
defparam \alu_b_mux_output[9]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N16
cycloneive_lcell_comb \alu_b_mux_output[8]~54 (
// Equation(s):
// alu_b_mux_output_8 = (\alu_b_mux_output[8]~53_combout ) # ((!always06 & (!forwardb_1 & temp_rdat_two_output_8)))

	.dataa(always04),
	.datab(\alu_b_mux_output[8]~53_combout ),
	.datac(forwardb_1),
	.datad(temp_rdat_two_output_8),
	.cin(gnd),
	.combout(alu_b_mux_output_8),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[8]~54 .lut_mask = 16'hCDCC;
defparam \alu_b_mux_output[8]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N20
cycloneive_lcell_comb \alu_b_mux_output[7]~56 (
// Equation(s):
// alu_b_mux_output_7 = (\alu_b_mux_output[7]~55_combout ) # ((!always06 & (temp_rdat_two_output_7 & !forwardb_1)))

	.dataa(always04),
	.datab(temp_rdat_two_output_7),
	.datac(forwardb_1),
	.datad(\alu_b_mux_output[7]~55_combout ),
	.cin(gnd),
	.combout(alu_b_mux_output_7),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[7]~56 .lut_mask = 16'hFF04;
defparam \alu_b_mux_output[7]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N22
cycloneive_lcell_comb \alu_b_mux_output[6]~58 (
// Equation(s):
// alu_b_mux_output_6 = (\alu_b_mux_output[6]~57_combout ) # ((!always06 & (!forwardb_1 & temp_rdat_two_output_6)))

	.dataa(\alu_b_mux_output[6]~57_combout ),
	.datab(always04),
	.datac(forwardb_1),
	.datad(temp_rdat_two_output_6),
	.cin(gnd),
	.combout(alu_b_mux_output_6),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[6]~58 .lut_mask = 16'hABAA;
defparam \alu_b_mux_output[6]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N6
cycloneive_lcell_comb \alu_b_mux_output[5]~60 (
// Equation(s):
// alu_b_mux_output_5 = (\alu_b_mux_output[5]~59_combout ) # ((temp_rdat_two_output_5 & (!always06 & !forwardb_1)))

	.dataa(\alu_b_mux_output[5]~59_combout ),
	.datab(temp_rdat_two_output_5),
	.datac(always04),
	.datad(forwardb_1),
	.cin(gnd),
	.combout(alu_b_mux_output_5),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[5]~60 .lut_mask = 16'hAAAE;
defparam \alu_b_mux_output[5]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N0
cycloneive_lcell_comb \alu_b_mux_output[13]~62 (
// Equation(s):
// alu_b_mux_output_13 = (\alu_b_mux_output[13]~61_combout ) # ((!forwardb_1 & (!always06 & temp_rdat_two_output_13)))

	.dataa(forwardb_1),
	.datab(\alu_b_mux_output[13]~61_combout ),
	.datac(always04),
	.datad(temp_rdat_two_output_13),
	.cin(gnd),
	.combout(alu_b_mux_output_13),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[13]~62 .lut_mask = 16'hCDCC;
defparam \alu_b_mux_output[13]~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N8
cycloneive_lcell_comb \alu_b_mux_output[11]~64 (
// Equation(s):
// alu_b_mux_output_111 = (\alu_b_mux_output[11]~63_combout ) # ((!always06 & (temp_rdat_two_output_11 & !forwardb_1)))

	.dataa(\alu_b_mux_output[11]~63_combout ),
	.datab(always04),
	.datac(temp_rdat_two_output_11),
	.datad(forwardb_1),
	.cin(gnd),
	.combout(alu_b_mux_output_111),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[11]~64 .lut_mask = 16'hAABA;
defparam \alu_b_mux_output[11]~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N0
cycloneive_lcell_comb \alu_b_mux_output[2]~4 (
// Equation(s):
// \alu_b_mux_output[2]~4_combout  = (forwardb_1 & (!always06 & (Mux29))) # (!forwardb_1 & (always06 & ((temp_aluResult_2))))

	.dataa(forwardb_1),
	.datab(always04),
	.datac(Mux29),
	.datad(temp_aluResult_2),
	.cin(gnd),
	.combout(\alu_b_mux_output[2]~4_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[2]~4 .lut_mask = 16'h6420;
defparam \alu_b_mux_output[2]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N4
cycloneive_lcell_comb \alu_b_mux_output[3]~6 (
// Equation(s):
// \alu_b_mux_output[3]~6_combout  = (forwardb_1 & (((Mux28 & !always06)))) # (!forwardb_1 & (temp_aluResult_3 & ((always06))))

	.dataa(temp_aluResult_3),
	.datab(Mux28),
	.datac(forwardb_1),
	.datad(always04),
	.cin(gnd),
	.combout(\alu_b_mux_output[3]~6_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[3]~6 .lut_mask = 16'h0AC0;
defparam \alu_b_mux_output[3]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N30
cycloneive_lcell_comb \alu_b_mux_output[4]~8 (
// Equation(s):
// \alu_b_mux_output[4]~8_combout  = (forwardb_1 & (((Mux27 & !always06)))) # (!forwardb_1 & (temp_aluResult_4 & ((always06))))

	.dataa(forwardb_1),
	.datab(temp_aluResult_4),
	.datac(Mux27),
	.datad(always04),
	.cin(gnd),
	.combout(\alu_b_mux_output[4]~8_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[4]~8 .lut_mask = 16'h44A0;
defparam \alu_b_mux_output[4]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N4
cycloneive_lcell_comb \alu_b_mux_output[15]~10 (
// Equation(s):
// \alu_b_mux_output[15]~10_combout  = (forwardb_1 & (!always06 & ((Mux16)))) # (!forwardb_1 & (always06 & (temp_aluResult_15)))

	.dataa(forwardb_1),
	.datab(always04),
	.datac(temp_aluResult_15),
	.datad(Mux16),
	.cin(gnd),
	.combout(\alu_b_mux_output[15]~10_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[15]~10 .lut_mask = 16'h6240;
defparam \alu_b_mux_output[15]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N12
cycloneive_lcell_comb \alu_b_mux_output[12]~12 (
// Equation(s):
// \alu_b_mux_output[12]~12_combout  = (always06 & (((temp_aluResult_12 & !forwardb_1)))) # (!always06 & (Mux19 & ((forwardb_1))))

	.dataa(Mux19),
	.datab(always04),
	.datac(temp_aluResult_12),
	.datad(forwardb_1),
	.cin(gnd),
	.combout(\alu_b_mux_output[12]~12_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[12]~12 .lut_mask = 16'h22C0;
defparam \alu_b_mux_output[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N8
cycloneive_lcell_comb \alu_b_mux_output[27]~14 (
// Equation(s):
// \alu_b_mux_output[27]~14_combout  = (always0) # ((!always06 & ((!always01) # (!always03))))

	.dataa(always04),
	.datab(always03),
	.datac(always01),
	.datad(always0),
	.cin(gnd),
	.combout(\alu_b_mux_output[27]~14_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[27]~14 .lut_mask = 16'hFF15;
defparam \alu_b_mux_output[27]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N6
cycloneive_lcell_comb \alu_b_mux_output[27]~15 (
// Equation(s):
// \alu_b_mux_output[27]~15_combout  = (forwardb_1 & ((Mux4) # ((\alu_b_mux_output[27]~14_combout )))) # (!forwardb_1 & (((temp_aluResult_27 & !\alu_b_mux_output[27]~14_combout ))))

	.dataa(Mux4),
	.datab(forwardb_1),
	.datac(temp_aluResult_27),
	.datad(\alu_b_mux_output[27]~14_combout ),
	.cin(gnd),
	.combout(\alu_b_mux_output[27]~15_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[27]~15 .lut_mask = 16'hCCB8;
defparam \alu_b_mux_output[27]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N18
cycloneive_lcell_comb \alu_b_mux_output[18]~17 (
// Equation(s):
// \alu_b_mux_output[18]~17_combout  = (\alu_b_mux_output[27]~14_combout  & (((forwardb_1)))) # (!\alu_b_mux_output[27]~14_combout  & ((forwardb_1 & (Mux13)) # (!forwardb_1 & ((temp_aluResult_18)))))

	.dataa(Mux13),
	.datab(temp_aluResult_18),
	.datac(\alu_b_mux_output[27]~14_combout ),
	.datad(forwardb_1),
	.cin(gnd),
	.combout(\alu_b_mux_output[18]~17_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[18]~17 .lut_mask = 16'hFA0C;
defparam \alu_b_mux_output[18]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N24
cycloneive_lcell_comb \alu_b_mux_output[17]~19 (
// Equation(s):
// \alu_b_mux_output[17]~19_combout  = (\alu_b_mux_output[27]~14_combout  & (((forwardb_1)))) # (!\alu_b_mux_output[27]~14_combout  & ((forwardb_1 & ((Mux14))) # (!forwardb_1 & (temp_aluResult_17))))

	.dataa(temp_aluResult_17),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(Mux14),
	.datad(forwardb_1),
	.cin(gnd),
	.combout(\alu_b_mux_output[17]~19_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[17]~19 .lut_mask = 16'hFC22;
defparam \alu_b_mux_output[17]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N4
cycloneive_lcell_comb \alu_b_mux_output[16]~21 (
// Equation(s):
// \alu_b_mux_output[16]~21_combout  = (forwardb_1 & (((Mux15) # (\alu_b_mux_output[27]~14_combout )))) # (!forwardb_1 & (temp_aluResult_16 & ((!\alu_b_mux_output[27]~14_combout ))))

	.dataa(forwardb_1),
	.datab(temp_aluResult_16),
	.datac(Mux15),
	.datad(\alu_b_mux_output[27]~14_combout ),
	.cin(gnd),
	.combout(\alu_b_mux_output[16]~21_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[16]~21 .lut_mask = 16'hAAE4;
defparam \alu_b_mux_output[16]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N14
cycloneive_lcell_comb \alu_b_mux_output[31]~23 (
// Equation(s):
// \alu_b_mux_output[31]~23_combout  = (forwardb_1 & ((\alu_b_mux_output[27]~14_combout ) # ((Mux0)))) # (!forwardb_1 & (!\alu_b_mux_output[27]~14_combout  & ((temp_aluResult_31))))

	.dataa(forwardb_1),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(Mux0),
	.datad(temp_aluResult_31),
	.cin(gnd),
	.combout(\alu_b_mux_output[31]~23_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[31]~23 .lut_mask = 16'hB9A8;
defparam \alu_b_mux_output[31]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N24
cycloneive_lcell_comb \alu_b_mux_output[30]~25 (
// Equation(s):
// \alu_b_mux_output[30]~25_combout  = (\alu_b_mux_output[27]~14_combout  & (((forwardb_1)))) # (!\alu_b_mux_output[27]~14_combout  & ((forwardb_1 & (Mux1)) # (!forwardb_1 & ((temp_aluResult_30)))))

	.dataa(Mux1),
	.datab(temp_aluResult_30),
	.datac(\alu_b_mux_output[27]~14_combout ),
	.datad(forwardb_1),
	.cin(gnd),
	.combout(\alu_b_mux_output[30]~25_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[30]~25 .lut_mask = 16'hFA0C;
defparam \alu_b_mux_output[30]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N30
cycloneive_lcell_comb \alu_b_mux_output[29]~27 (
// Equation(s):
// \alu_b_mux_output[29]~27_combout  = (forwardb_1 & ((Mux2) # ((\alu_b_mux_output[27]~14_combout )))) # (!forwardb_1 & (((!\alu_b_mux_output[27]~14_combout  & temp_aluResult_29))))

	.dataa(Mux2),
	.datab(forwardb_1),
	.datac(\alu_b_mux_output[27]~14_combout ),
	.datad(temp_aluResult_29),
	.cin(gnd),
	.combout(\alu_b_mux_output[29]~27_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[29]~27 .lut_mask = 16'hCBC8;
defparam \alu_b_mux_output[29]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N6
cycloneive_lcell_comb \alu_b_mux_output[28]~29 (
// Equation(s):
// \alu_b_mux_output[28]~29_combout  = (forwardb_1 & ((\alu_b_mux_output[27]~14_combout ) # ((Mux3)))) # (!forwardb_1 & (!\alu_b_mux_output[27]~14_combout  & ((temp_aluResult_28))))

	.dataa(forwardb_1),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(Mux3),
	.datad(temp_aluResult_28),
	.cin(gnd),
	.combout(\alu_b_mux_output[28]~29_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[28]~29 .lut_mask = 16'hB9A8;
defparam \alu_b_mux_output[28]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N26
cycloneive_lcell_comb \alu_b_mux_output[26]~31 (
// Equation(s):
// \alu_b_mux_output[26]~31_combout  = (forwardb_1 & ((\alu_b_mux_output[27]~14_combout ) # ((Mux5)))) # (!forwardb_1 & (!\alu_b_mux_output[27]~14_combout  & (temp_aluResult_26)))

	.dataa(forwardb_1),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(temp_aluResult_26),
	.datad(Mux5),
	.cin(gnd),
	.combout(\alu_b_mux_output[26]~31_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[26]~31 .lut_mask = 16'hBA98;
defparam \alu_b_mux_output[26]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N14
cycloneive_lcell_comb \alu_b_mux_output[25]~33 (
// Equation(s):
// \alu_b_mux_output[25]~33_combout  = (forwardb_1 & ((Mux6) # ((\alu_b_mux_output[27]~14_combout )))) # (!forwardb_1 & (((temp_aluResult_25 & !\alu_b_mux_output[27]~14_combout ))))

	.dataa(Mux6),
	.datab(temp_aluResult_25),
	.datac(forwardb_1),
	.datad(\alu_b_mux_output[27]~14_combout ),
	.cin(gnd),
	.combout(\alu_b_mux_output[25]~33_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[25]~33 .lut_mask = 16'hF0AC;
defparam \alu_b_mux_output[25]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N10
cycloneive_lcell_comb \alu_b_mux_output[24]~35 (
// Equation(s):
// \alu_b_mux_output[24]~35_combout  = (\alu_b_mux_output[27]~14_combout  & (forwardb_1)) # (!\alu_b_mux_output[27]~14_combout  & ((forwardb_1 & ((Mux7))) # (!forwardb_1 & (temp_aluResult_24))))

	.dataa(\alu_b_mux_output[27]~14_combout ),
	.datab(forwardb_1),
	.datac(temp_aluResult_24),
	.datad(Mux7),
	.cin(gnd),
	.combout(\alu_b_mux_output[24]~35_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[24]~35 .lut_mask = 16'hDC98;
defparam \alu_b_mux_output[24]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N10
cycloneive_lcell_comb \alu_b_mux_output[23]~37 (
// Equation(s):
// \alu_b_mux_output[23]~37_combout  = (forwardb_1 & ((\alu_b_mux_output[27]~14_combout ) # ((Mux8)))) # (!forwardb_1 & (!\alu_b_mux_output[27]~14_combout  & (temp_aluResult_23)))

	.dataa(forwardb_1),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(temp_aluResult_23),
	.datad(Mux8),
	.cin(gnd),
	.combout(\alu_b_mux_output[23]~37_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[23]~37 .lut_mask = 16'hBA98;
defparam \alu_b_mux_output[23]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N8
cycloneive_lcell_comb \alu_b_mux_output[22]~39 (
// Equation(s):
// \alu_b_mux_output[22]~39_combout  = (forwardb_1 & ((\alu_b_mux_output[27]~14_combout ) # ((Mux9)))) # (!forwardb_1 & (!\alu_b_mux_output[27]~14_combout  & ((temp_aluResult_22))))

	.dataa(forwardb_1),
	.datab(\alu_b_mux_output[27]~14_combout ),
	.datac(Mux9),
	.datad(temp_aluResult_22),
	.cin(gnd),
	.combout(\alu_b_mux_output[22]~39_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[22]~39 .lut_mask = 16'hB9A8;
defparam \alu_b_mux_output[22]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N18
cycloneive_lcell_comb \alu_b_mux_output[21]~41 (
// Equation(s):
// \alu_b_mux_output[21]~41_combout  = (\alu_b_mux_output[27]~14_combout  & (((forwardb_1)))) # (!\alu_b_mux_output[27]~14_combout  & ((forwardb_1 & ((Mux10))) # (!forwardb_1 & (temp_aluResult_21))))

	.dataa(\alu_b_mux_output[27]~14_combout ),
	.datab(temp_aluResult_21),
	.datac(Mux10),
	.datad(forwardb_1),
	.cin(gnd),
	.combout(\alu_b_mux_output[21]~41_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[21]~41 .lut_mask = 16'hFA44;
defparam \alu_b_mux_output[21]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N6
cycloneive_lcell_comb \alu_b_mux_output[20]~43 (
// Equation(s):
// \alu_b_mux_output[20]~43_combout  = (forwardb_1 & ((Mux11) # ((\alu_b_mux_output[27]~14_combout )))) # (!forwardb_1 & (((!\alu_b_mux_output[27]~14_combout  & temp_aluResult_20))))

	.dataa(Mux11),
	.datab(forwardb_1),
	.datac(\alu_b_mux_output[27]~14_combout ),
	.datad(temp_aluResult_20),
	.cin(gnd),
	.combout(\alu_b_mux_output[20]~43_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[20]~43 .lut_mask = 16'hCBC8;
defparam \alu_b_mux_output[20]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N22
cycloneive_lcell_comb \alu_b_mux_output[19]~45 (
// Equation(s):
// \alu_b_mux_output[19]~45_combout  = (forwardb_1 & ((Mux12) # ((\alu_b_mux_output[27]~14_combout )))) # (!forwardb_1 & (((temp_aluResult_19 & !\alu_b_mux_output[27]~14_combout ))))

	.dataa(Mux12),
	.datab(temp_aluResult_19),
	.datac(forwardb_1),
	.datad(\alu_b_mux_output[27]~14_combout ),
	.cin(gnd),
	.combout(\alu_b_mux_output[19]~45_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[19]~45 .lut_mask = 16'hF0AC;
defparam \alu_b_mux_output[19]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N22
cycloneive_lcell_comb \alu_b_mux_output[10]~47 (
// Equation(s):
// \alu_b_mux_output[10]~47_combout  = (forwardb_1 & (Mux21 & ((!always06)))) # (!forwardb_1 & (((temp_aluResult_10 & always06))))

	.dataa(forwardb_1),
	.datab(Mux21),
	.datac(temp_aluResult_10),
	.datad(always04),
	.cin(gnd),
	.combout(\alu_b_mux_output[10]~47_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[10]~47 .lut_mask = 16'h5088;
defparam \alu_b_mux_output[10]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N10
cycloneive_lcell_comb \alu_b_mux_output[14]~49 (
// Equation(s):
// \alu_b_mux_output[14]~49_combout  = (always06 & (temp_aluResult_14 & (!forwardb_1))) # (!always06 & (((forwardb_1 & Mux17))))

	.dataa(temp_aluResult_14),
	.datab(always04),
	.datac(forwardb_1),
	.datad(Mux17),
	.cin(gnd),
	.combout(\alu_b_mux_output[14]~49_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[14]~49 .lut_mask = 16'h3808;
defparam \alu_b_mux_output[14]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N2
cycloneive_lcell_comb \alu_b_mux_output[9]~51 (
// Equation(s):
// \alu_b_mux_output[9]~51_combout  = (always06 & (temp_aluResult_9 & (!forwardb_1))) # (!always06 & (((forwardb_1 & Mux22))))

	.dataa(always04),
	.datab(temp_aluResult_9),
	.datac(forwardb_1),
	.datad(Mux22),
	.cin(gnd),
	.combout(\alu_b_mux_output[9]~51_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[9]~51 .lut_mask = 16'h5808;
defparam \alu_b_mux_output[9]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N20
cycloneive_lcell_comb \alu_b_mux_output[8]~53 (
// Equation(s):
// \alu_b_mux_output[8]~53_combout  = (always06 & (((!forwardb_1 & temp_aluResult_8)))) # (!always06 & (Mux23 & (forwardb_1)))

	.dataa(always04),
	.datab(Mux23),
	.datac(forwardb_1),
	.datad(temp_aluResult_8),
	.cin(gnd),
	.combout(\alu_b_mux_output[8]~53_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[8]~53 .lut_mask = 16'h4A40;
defparam \alu_b_mux_output[8]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N0
cycloneive_lcell_comb \alu_b_mux_output[7]~55 (
// Equation(s):
// \alu_b_mux_output[7]~55_combout  = (always06 & (temp_aluResult_7 & (!forwardb_1))) # (!always06 & (((forwardb_1 & Mux24))))

	.dataa(always04),
	.datab(temp_aluResult_7),
	.datac(forwardb_1),
	.datad(Mux24),
	.cin(gnd),
	.combout(\alu_b_mux_output[7]~55_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[7]~55 .lut_mask = 16'h5808;
defparam \alu_b_mux_output[7]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N6
cycloneive_lcell_comb \alu_b_mux_output[6]~57 (
// Equation(s):
// \alu_b_mux_output[6]~57_combout  = (forwardb_1 & (((!always06 & Mux25)))) # (!forwardb_1 & (temp_aluResult_6 & (always06)))

	.dataa(forwardb_1),
	.datab(temp_aluResult_6),
	.datac(always04),
	.datad(Mux25),
	.cin(gnd),
	.combout(\alu_b_mux_output[6]~57_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[6]~57 .lut_mask = 16'h4A40;
defparam \alu_b_mux_output[6]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N22
cycloneive_lcell_comb \alu_b_mux_output[5]~59 (
// Equation(s):
// \alu_b_mux_output[5]~59_combout  = (always06 & (temp_aluResult_5 & ((!forwardb_1)))) # (!always06 & (((Mux26 & forwardb_1))))

	.dataa(always04),
	.datab(temp_aluResult_5),
	.datac(Mux26),
	.datad(forwardb_1),
	.cin(gnd),
	.combout(\alu_b_mux_output[5]~59_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[5]~59 .lut_mask = 16'h5088;
defparam \alu_b_mux_output[5]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N28
cycloneive_lcell_comb \alu_b_mux_output[13]~61 (
// Equation(s):
// \alu_b_mux_output[13]~61_combout  = (forwardb_1 & (!always06 & ((Mux18)))) # (!forwardb_1 & (always06 & (temp_aluResult_13)))

	.dataa(forwardb_1),
	.datab(always04),
	.datac(temp_aluResult_13),
	.datad(Mux18),
	.cin(gnd),
	.combout(\alu_b_mux_output[13]~61_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[13]~61 .lut_mask = 16'h6240;
defparam \alu_b_mux_output[13]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N12
cycloneive_lcell_comb \alu_b_mux_output[11]~63 (
// Equation(s):
// \alu_b_mux_output[11]~63_combout  = (always06 & (((temp_aluResult_11 & !forwardb_1)))) # (!always06 & (Mux20 & ((forwardb_1))))

	.dataa(Mux20),
	.datab(always04),
	.datac(temp_aluResult_11),
	.datad(forwardb_1),
	.cin(gnd),
	.combout(\alu_b_mux_output[11]~63_combout ),
	.cout());
// synopsys translate_off
defparam \alu_b_mux_output[11]~63 .lut_mask = 16'h22C0;
defparam \alu_b_mux_output[11]~63 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module alu_source_mux (
	temp_signzerovalue_output_16,
	temp_imemload_output_1,
	temp_imemload_output_7,
	temp_ALUsrc_output_1,
	temp_ALUsrc_output_0,
	Mux30,
	alu_b_mux_output_1,
	alu_b_mux_output_11,
	Mux16,
	Mux301,
	alu_b_mux_output_0,
	temp_imemload_output_0,
	temp_imemload_output_6,
	Mux31,
	alu_b_mux_output_01,
	Mux311,
	temp_imemload_output_2,
	temp_imemload_output_8,
	Mux29,
	alu_b_mux_output_2,
	Mux291,
	temp_imemload_output_3,
	temp_imemload_output_9,
	Mux28,
	alu_b_mux_output_3,
	Mux281,
	temp_imemload_output_4,
	temp_imemload_output_10,
	Mux27,
	alu_b_mux_output_4,
	Mux271,
	alu_b_mux_output_15,
	temp_imemload_output_15,
	Mux161,
	alu_b_mux_output_12,
	temp_imemload_output_12,
	Mux19,
	alu_b_mux_output_27,
	Mux4,
	alu_b_mux_output_18,
	Mux13,
	alu_b_mux_output_17,
	Mux14,
	alu_b_mux_output_16,
	Mux15,
	alu_b_mux_output_31,
	Mux0,
	alu_b_mux_output_30,
	Mux1,
	alu_b_mux_output_29,
	Mux2,
	alu_b_mux_output_28,
	Mux3,
	alu_b_mux_output_26,
	Mux5,
	alu_b_mux_output_25,
	Mux6,
	alu_b_mux_output_24,
	Mux7,
	alu_b_mux_output_23,
	Mux8,
	alu_b_mux_output_22,
	Mux9,
	alu_b_mux_output_21,
	Mux10,
	alu_b_mux_output_20,
	Mux11,
	alu_b_mux_output_19,
	Mux12,
	temp_imemload_output_14,
	Mux17,
	alu_b_mux_output_10,
	Mux21,
	alu_b_mux_output_14,
	alu_b_mux_output_9,
	Mux22,
	alu_b_mux_output_8,
	Mux23,
	alu_b_mux_output_7,
	Mux24,
	alu_b_mux_output_6,
	Mux25,
	alu_b_mux_output_5,
	temp_imemload_output_5,
	Mux26,
	alu_b_mux_output_13,
	temp_imemload_output_13,
	Mux18,
	alu_b_mux_output_111,
	temp_imemload_output_11,
	Mux20,
	Mux171,
	devpor,
	devclrn,
	devoe);
input 	temp_signzerovalue_output_16;
input 	temp_imemload_output_1;
input 	temp_imemload_output_7;
input 	temp_ALUsrc_output_1;
input 	temp_ALUsrc_output_0;
output 	Mux30;
input 	alu_b_mux_output_1;
input 	alu_b_mux_output_11;
output 	Mux16;
output 	Mux301;
input 	alu_b_mux_output_0;
input 	temp_imemload_output_0;
input 	temp_imemload_output_6;
output 	Mux31;
input 	alu_b_mux_output_01;
output 	Mux311;
input 	temp_imemload_output_2;
input 	temp_imemload_output_8;
output 	Mux29;
input 	alu_b_mux_output_2;
output 	Mux291;
input 	temp_imemload_output_3;
input 	temp_imemload_output_9;
output 	Mux28;
input 	alu_b_mux_output_3;
output 	Mux281;
input 	temp_imemload_output_4;
input 	temp_imemload_output_10;
output 	Mux27;
input 	alu_b_mux_output_4;
output 	Mux271;
input 	alu_b_mux_output_15;
input 	temp_imemload_output_15;
output 	Mux161;
input 	alu_b_mux_output_12;
input 	temp_imemload_output_12;
output 	Mux19;
input 	alu_b_mux_output_27;
output 	Mux4;
input 	alu_b_mux_output_18;
output 	Mux13;
input 	alu_b_mux_output_17;
output 	Mux14;
input 	alu_b_mux_output_16;
output 	Mux15;
input 	alu_b_mux_output_31;
output 	Mux0;
input 	alu_b_mux_output_30;
output 	Mux1;
input 	alu_b_mux_output_29;
output 	Mux2;
input 	alu_b_mux_output_28;
output 	Mux3;
input 	alu_b_mux_output_26;
output 	Mux5;
input 	alu_b_mux_output_25;
output 	Mux6;
input 	alu_b_mux_output_24;
output 	Mux7;
input 	alu_b_mux_output_23;
output 	Mux8;
input 	alu_b_mux_output_22;
output 	Mux9;
input 	alu_b_mux_output_21;
output 	Mux10;
input 	alu_b_mux_output_20;
output 	Mux11;
input 	alu_b_mux_output_19;
output 	Mux12;
input 	temp_imemload_output_14;
output 	Mux17;
input 	alu_b_mux_output_10;
output 	Mux21;
input 	alu_b_mux_output_14;
input 	alu_b_mux_output_9;
output 	Mux22;
input 	alu_b_mux_output_8;
output 	Mux23;
input 	alu_b_mux_output_7;
output 	Mux24;
input 	alu_b_mux_output_6;
output 	Mux25;
input 	alu_b_mux_output_5;
input 	temp_imemload_output_5;
output 	Mux26;
input 	alu_b_mux_output_13;
input 	temp_imemload_output_13;
output 	Mux18;
input 	alu_b_mux_output_111;
input 	temp_imemload_output_11;
output 	Mux20;
output 	Mux171;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X61_Y39_N26
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// Mux30 = (temp_ALUsrc_output_1 & (!temp_ALUsrc_output_0 & (temp_imemload_output_7))) # (!temp_ALUsrc_output_1 & (temp_ALUsrc_output_0 & ((temp_imemload_output_1))))

	.dataa(temp_ALUsrc_output_1),
	.datab(temp_ALUsrc_output_0),
	.datac(temp_imemload_output_7),
	.datad(temp_imemload_output_1),
	.cin(gnd),
	.combout(Mux30),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'h6420;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N14
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// Mux16 = temp_ALUsrc_output_1 $ (temp_ALUsrc_output_0)

	.dataa(temp_ALUsrc_output_1),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_ALUsrc_output_0),
	.cin(gnd),
	.combout(Mux16),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'h55AA;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N10
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// Mux301 = (Mux30) # ((!Mux16 & ((alu_b_mux_output_11) # (alu_b_mux_output_1))))

	.dataa(Mux16),
	.datab(alu_b_mux_output_11),
	.datac(Mux30),
	.datad(alu_b_mux_output_1),
	.cin(gnd),
	.combout(Mux301),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hF5F4;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N12
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// Mux31 = (temp_ALUsrc_output_1 & (((temp_imemload_output_6 & !temp_ALUsrc_output_0)))) # (!temp_ALUsrc_output_1 & (temp_imemload_output_0 & ((temp_ALUsrc_output_0))))

	.dataa(temp_ALUsrc_output_1),
	.datab(temp_imemload_output_0),
	.datac(temp_imemload_output_6),
	.datad(temp_ALUsrc_output_0),
	.cin(gnd),
	.combout(Mux31),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'h44A0;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N14
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// Mux311 = (Mux31) # ((!Mux16 & ((alu_b_mux_output_01) # (alu_b_mux_output_0))))

	.dataa(Mux31),
	.datab(alu_b_mux_output_01),
	.datac(alu_b_mux_output_0),
	.datad(Mux16),
	.cin(gnd),
	.combout(Mux311),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hAAFE;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N26
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// Mux29 = (temp_ALUsrc_output_1 & (((temp_imemload_output_8 & !temp_ALUsrc_output_0)))) # (!temp_ALUsrc_output_1 & (temp_imemload_output_2 & ((temp_ALUsrc_output_0))))

	.dataa(temp_imemload_output_2),
	.datab(temp_imemload_output_8),
	.datac(temp_ALUsrc_output_1),
	.datad(temp_ALUsrc_output_0),
	.cin(gnd),
	.combout(Mux29),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'h0AC0;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N20
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// Mux291 = (Mux29) # ((alu_b_mux_output_2 & (temp_ALUsrc_output_0 $ (!temp_ALUsrc_output_1))))

	.dataa(Mux29),
	.datab(temp_ALUsrc_output_0),
	.datac(temp_ALUsrc_output_1),
	.datad(alu_b_mux_output_2),
	.cin(gnd),
	.combout(Mux291),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hEBAA;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N30
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// Mux28 = (temp_ALUsrc_output_1 & (((temp_imemload_output_9 & !temp_ALUsrc_output_0)))) # (!temp_ALUsrc_output_1 & (temp_imemload_output_3 & ((temp_ALUsrc_output_0))))

	.dataa(temp_imemload_output_3),
	.datab(temp_imemload_output_9),
	.datac(temp_ALUsrc_output_1),
	.datad(temp_ALUsrc_output_0),
	.cin(gnd),
	.combout(Mux28),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'h0AC0;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N12
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// Mux281 = (Mux28) # ((alu_b_mux_output_3 & (temp_ALUsrc_output_0 $ (!temp_ALUsrc_output_1))))

	.dataa(Mux28),
	.datab(temp_ALUsrc_output_0),
	.datac(temp_ALUsrc_output_1),
	.datad(alu_b_mux_output_3),
	.cin(gnd),
	.combout(Mux281),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hEBAA;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N26
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// Mux27 = (temp_ALUsrc_output_0 & (((!temp_ALUsrc_output_1 & temp_imemload_output_4)))) # (!temp_ALUsrc_output_0 & (temp_imemload_output_10 & (temp_ALUsrc_output_1)))

	.dataa(temp_imemload_output_10),
	.datab(temp_ALUsrc_output_0),
	.datac(temp_ALUsrc_output_1),
	.datad(temp_imemload_output_4),
	.cin(gnd),
	.combout(Mux27),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'h2C20;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N8
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// Mux271 = (Mux27) # ((alu_b_mux_output_4 & (temp_ALUsrc_output_0 $ (!temp_ALUsrc_output_1))))

	.dataa(temp_ALUsrc_output_0),
	.datab(temp_ALUsrc_output_1),
	.datac(Mux27),
	.datad(alu_b_mux_output_4),
	.cin(gnd),
	.combout(Mux271),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hF9F0;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N14
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// Mux161 = (temp_ALUsrc_output_1 & (((temp_ALUsrc_output_0 & alu_b_mux_output_15)))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & (temp_imemload_output_15)) # (!temp_ALUsrc_output_0 & ((alu_b_mux_output_15)))))

	.dataa(temp_ALUsrc_output_1),
	.datab(temp_imemload_output_15),
	.datac(temp_ALUsrc_output_0),
	.datad(alu_b_mux_output_15),
	.cin(gnd),
	.combout(Mux161),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hE540;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N16
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// Mux19 = (temp_ALUsrc_output_1 & (((temp_ALUsrc_output_0 & alu_b_mux_output_12)))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & (temp_imemload_output_12)) # (!temp_ALUsrc_output_0 & ((alu_b_mux_output_12)))))

	.dataa(temp_ALUsrc_output_1),
	.datab(temp_imemload_output_12),
	.datac(temp_ALUsrc_output_0),
	.datad(alu_b_mux_output_12),
	.cin(gnd),
	.combout(Mux19),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hE540;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N12
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// Mux4 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & ((alu_b_mux_output_27))) # (!temp_ALUsrc_output_1 & (temp_signzerovalue_output_16)))) # (!temp_ALUsrc_output_0 & (((alu_b_mux_output_27 & !temp_ALUsrc_output_1))))

	.dataa(temp_ALUsrc_output_0),
	.datab(temp_signzerovalue_output_16),
	.datac(alu_b_mux_output_27),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux4),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hA0D8;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N10
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// Mux13 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & (alu_b_mux_output_18)) # (!temp_ALUsrc_output_1 & ((temp_signzerovalue_output_16))))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_18 & ((!temp_ALUsrc_output_1))))

	.dataa(temp_ALUsrc_output_0),
	.datab(alu_b_mux_output_18),
	.datac(temp_signzerovalue_output_16),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux13),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'h88E4;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N16
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// Mux14 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & ((alu_b_mux_output_17))) # (!temp_ALUsrc_output_1 & (temp_signzerovalue_output_16)))) # (!temp_ALUsrc_output_0 & (((alu_b_mux_output_17 & !temp_ALUsrc_output_1))))

	.dataa(temp_ALUsrc_output_0),
	.datab(temp_signzerovalue_output_16),
	.datac(alu_b_mux_output_17),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux14),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hA0D8;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N28
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// Mux15 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & ((alu_b_mux_output_16))) # (!temp_ALUsrc_output_1 & (temp_signzerovalue_output_16)))) # (!temp_ALUsrc_output_0 & (((!temp_ALUsrc_output_1 & alu_b_mux_output_16))))

	.dataa(temp_signzerovalue_output_16),
	.datab(temp_ALUsrc_output_0),
	.datac(temp_ALUsrc_output_1),
	.datad(alu_b_mux_output_16),
	.cin(gnd),
	.combout(Mux15),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hCB08;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N4
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// Mux0 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & (alu_b_mux_output_31)) # (!temp_ALUsrc_output_1 & ((temp_signzerovalue_output_16))))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_31 & ((!temp_ALUsrc_output_1))))

	.dataa(alu_b_mux_output_31),
	.datab(temp_signzerovalue_output_16),
	.datac(temp_ALUsrc_output_0),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux0),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hA0CA;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N4
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// Mux1 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & (alu_b_mux_output_30)) # (!temp_ALUsrc_output_1 & ((temp_signzerovalue_output_16))))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_30 & ((!temp_ALUsrc_output_1))))

	.dataa(temp_ALUsrc_output_0),
	.datab(alu_b_mux_output_30),
	.datac(temp_signzerovalue_output_16),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux1),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'h88E4;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N6
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// Mux2 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & (alu_b_mux_output_29)) # (!temp_ALUsrc_output_1 & ((temp_signzerovalue_output_16))))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_29 & ((!temp_ALUsrc_output_1))))

	.dataa(temp_ALUsrc_output_0),
	.datab(alu_b_mux_output_29),
	.datac(temp_signzerovalue_output_16),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux2),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'h88E4;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N22
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// Mux3 = (temp_ALUsrc_output_1 & (alu_b_mux_output_28 & (temp_ALUsrc_output_0))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & ((temp_signzerovalue_output_16))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_28))))

	.dataa(temp_ALUsrc_output_1),
	.datab(alu_b_mux_output_28),
	.datac(temp_ALUsrc_output_0),
	.datad(temp_signzerovalue_output_16),
	.cin(gnd),
	.combout(Mux3),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hD484;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N10
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// Mux5 = (temp_ALUsrc_output_1 & (alu_b_mux_output_26 & (temp_ALUsrc_output_0))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & ((temp_signzerovalue_output_16))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_26))))

	.dataa(temp_ALUsrc_output_1),
	.datab(alu_b_mux_output_26),
	.datac(temp_ALUsrc_output_0),
	.datad(temp_signzerovalue_output_16),
	.cin(gnd),
	.combout(Mux5),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hD484;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N26
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// Mux6 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & (alu_b_mux_output_25)) # (!temp_ALUsrc_output_1 & ((temp_signzerovalue_output_16))))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_25 & (!temp_ALUsrc_output_1)))

	.dataa(temp_ALUsrc_output_0),
	.datab(alu_b_mux_output_25),
	.datac(temp_ALUsrc_output_1),
	.datad(temp_signzerovalue_output_16),
	.cin(gnd),
	.combout(Mux6),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'h8E84;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N12
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// Mux7 = (temp_ALUsrc_output_1 & (((temp_ALUsrc_output_0 & alu_b_mux_output_24)))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & (temp_signzerovalue_output_16)) # (!temp_ALUsrc_output_0 & ((alu_b_mux_output_24)))))

	.dataa(temp_ALUsrc_output_1),
	.datab(temp_signzerovalue_output_16),
	.datac(temp_ALUsrc_output_0),
	.datad(alu_b_mux_output_24),
	.cin(gnd),
	.combout(Mux7),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hE540;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N26
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// Mux8 = (temp_ALUsrc_output_1 & (((alu_b_mux_output_23 & temp_ALUsrc_output_0)))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & (temp_signzerovalue_output_16)) # (!temp_ALUsrc_output_0 & ((alu_b_mux_output_23)))))

	.dataa(temp_signzerovalue_output_16),
	.datab(temp_ALUsrc_output_1),
	.datac(alu_b_mux_output_23),
	.datad(temp_ALUsrc_output_0),
	.cin(gnd),
	.combout(Mux8),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hE230;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N0
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// Mux9 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & (alu_b_mux_output_22)) # (!temp_ALUsrc_output_1 & ((temp_signzerovalue_output_16))))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_22 & ((!temp_ALUsrc_output_1))))

	.dataa(temp_ALUsrc_output_0),
	.datab(alu_b_mux_output_22),
	.datac(temp_signzerovalue_output_16),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux9),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'h88E4;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N28
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// Mux10 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & ((alu_b_mux_output_21))) # (!temp_ALUsrc_output_1 & (temp_signzerovalue_output_16)))) # (!temp_ALUsrc_output_0 & (((alu_b_mux_output_21 & !temp_ALUsrc_output_1))))

	.dataa(temp_signzerovalue_output_16),
	.datab(alu_b_mux_output_21),
	.datac(temp_ALUsrc_output_0),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux10),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hC0AC;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N14
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// Mux11 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & ((alu_b_mux_output_20))) # (!temp_ALUsrc_output_1 & (temp_signzerovalue_output_16)))) # (!temp_ALUsrc_output_0 & (((alu_b_mux_output_20 & !temp_ALUsrc_output_1))))

	.dataa(temp_signzerovalue_output_16),
	.datab(alu_b_mux_output_20),
	.datac(temp_ALUsrc_output_0),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux11),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hC0AC;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N20
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// Mux12 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & ((alu_b_mux_output_19))) # (!temp_ALUsrc_output_1 & (temp_signzerovalue_output_16)))) # (!temp_ALUsrc_output_0 & (((alu_b_mux_output_19 & !temp_ALUsrc_output_1))))

	.dataa(temp_signzerovalue_output_16),
	.datab(alu_b_mux_output_19),
	.datac(temp_ALUsrc_output_0),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux12),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hC0AC;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N24
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// Mux17 = (!temp_ALUsrc_output_1 & (temp_ALUsrc_output_0 & temp_imemload_output_14))

	.dataa(temp_ALUsrc_output_1),
	.datab(temp_ALUsrc_output_0),
	.datac(gnd),
	.datad(temp_imemload_output_14),
	.cin(gnd),
	.combout(Mux17),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'h4400;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N10
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// Mux21 = (temp_ALUsrc_output_1 & (alu_b_mux_output_10 & ((temp_ALUsrc_output_0)))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & ((temp_imemload_output_10))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_10))))

	.dataa(alu_b_mux_output_10),
	.datab(temp_ALUsrc_output_1),
	.datac(temp_imemload_output_10),
	.datad(temp_ALUsrc_output_0),
	.cin(gnd),
	.combout(Mux21),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hB822;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N16
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// Mux22 = (temp_ALUsrc_output_1 & (alu_b_mux_output_9 & (temp_ALUsrc_output_0))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & ((temp_imemload_output_9))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_9))))

	.dataa(alu_b_mux_output_9),
	.datab(temp_ALUsrc_output_1),
	.datac(temp_ALUsrc_output_0),
	.datad(temp_imemload_output_9),
	.cin(gnd),
	.combout(Mux22),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hB282;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N14
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// Mux23 = (temp_ALUsrc_output_1 & (alu_b_mux_output_8 & ((temp_ALUsrc_output_0)))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & ((temp_imemload_output_8))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_8))))

	.dataa(alu_b_mux_output_8),
	.datab(temp_imemload_output_8),
	.datac(temp_ALUsrc_output_1),
	.datad(temp_ALUsrc_output_0),
	.cin(gnd),
	.combout(Mux23),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hAC0A;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N16
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// Mux24 = (temp_ALUsrc_output_1 & (temp_ALUsrc_output_0 & ((alu_b_mux_output_7)))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & (temp_imemload_output_7)) # (!temp_ALUsrc_output_0 & ((alu_b_mux_output_7)))))

	.dataa(temp_ALUsrc_output_1),
	.datab(temp_ALUsrc_output_0),
	.datac(temp_imemload_output_7),
	.datad(alu_b_mux_output_7),
	.cin(gnd),
	.combout(Mux24),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hD940;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N20
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// Mux25 = (temp_ALUsrc_output_1 & (((alu_b_mux_output_6 & temp_ALUsrc_output_0)))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & (temp_imemload_output_6)) # (!temp_ALUsrc_output_0 & ((alu_b_mux_output_6)))))

	.dataa(temp_ALUsrc_output_1),
	.datab(temp_imemload_output_6),
	.datac(alu_b_mux_output_6),
	.datad(temp_ALUsrc_output_0),
	.cin(gnd),
	.combout(Mux25),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hE450;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N24
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// Mux26 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & (alu_b_mux_output_5)) # (!temp_ALUsrc_output_1 & ((temp_imemload_output_5))))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_5 & ((!temp_ALUsrc_output_1))))

	.dataa(alu_b_mux_output_5),
	.datab(temp_imemload_output_5),
	.datac(temp_ALUsrc_output_0),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux26),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hA0CA;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N30
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// Mux18 = (temp_ALUsrc_output_1 & (temp_ALUsrc_output_0 & ((alu_b_mux_output_13)))) # (!temp_ALUsrc_output_1 & ((temp_ALUsrc_output_0 & (temp_imemload_output_13)) # (!temp_ALUsrc_output_0 & ((alu_b_mux_output_13)))))

	.dataa(temp_ALUsrc_output_1),
	.datab(temp_ALUsrc_output_0),
	.datac(temp_imemload_output_13),
	.datad(alu_b_mux_output_13),
	.cin(gnd),
	.combout(Mux18),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hD940;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N30
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// Mux20 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & (alu_b_mux_output_111)) # (!temp_ALUsrc_output_1 & ((temp_imemload_output_11))))) # (!temp_ALUsrc_output_0 & (alu_b_mux_output_111 & ((!temp_ALUsrc_output_1))))

	.dataa(temp_ALUsrc_output_0),
	.datab(alu_b_mux_output_111),
	.datac(temp_imemload_output_11),
	.datad(temp_ALUsrc_output_1),
	.cin(gnd),
	.combout(Mux20),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'h88E4;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N6
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// Mux171 = (temp_ALUsrc_output_0 & ((temp_ALUsrc_output_1 & (alu_b_mux_output_14)) # (!temp_ALUsrc_output_1 & ((temp_imemload_output_14))))) # (!temp_ALUsrc_output_0 & (!temp_ALUsrc_output_1 & (alu_b_mux_output_14)))

	.dataa(temp_ALUsrc_output_0),
	.datab(temp_ALUsrc_output_1),
	.datac(alu_b_mux_output_14),
	.datad(temp_imemload_output_14),
	.cin(gnd),
	.combout(Mux171),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hB290;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module control_unit (
	temp_imemload_output_17,
	temp_imemload_output_16,
	temp_imemload_output_19,
	temp_imemload_output_18,
	temp_imemload_output_20,
	temp_imemload_output_22,
	temp_imemload_output_21,
	temp_imemload_output_24,
	temp_imemload_output_23,
	temp_imemload_output_25,
	temp_imemload_output_29,
	temp_imemload_output_31,
	temp_imemload_output_30,
	temp_imemload_output_28,
	Equal3,
	temp_imemload_output_27,
	temp_imemload_output_26,
	temp_branch_output,
	temp_imemload_output_0,
	temp_imemload_output_2,
	temp_imemload_output_3,
	temp_imemload_output_5,
	Equal31,
	temp_imemload_output_15,
	temp_imemload_output_14,
	temp_imemload_output_13,
	temp_imemload_output_12,
	temp_imemload_output_11,
	temp_imemload_output_10,
	temp_imemload_output_9,
	temp_imemload_output_8,
	temp_imemload_output_7,
	temp_imemload_output_6,
	temp_imemload_output_1,
	temp_imemload_output_4,
	Equal32,
	WideOr8,
	WideOr2,
	WideOr4,
	WideOr7,
	WideOr1,
	WideOr5,
	WideOr6,
	WideOr0,
	halt_out,
	halt_out1,
	WideOr3,
	WideOr10,
	memtoreg,
	WideOr9,
	devpor,
	devclrn,
	devoe);
input 	temp_imemload_output_17;
input 	temp_imemload_output_16;
input 	temp_imemload_output_19;
input 	temp_imemload_output_18;
input 	temp_imemload_output_20;
input 	temp_imemload_output_22;
input 	temp_imemload_output_21;
input 	temp_imemload_output_24;
input 	temp_imemload_output_23;
input 	temp_imemload_output_25;
input 	temp_imemload_output_29;
input 	temp_imemload_output_31;
input 	temp_imemload_output_30;
input 	temp_imemload_output_28;
output 	Equal3;
input 	temp_imemload_output_27;
input 	temp_imemload_output_26;
input 	temp_branch_output;
input 	temp_imemload_output_0;
input 	temp_imemload_output_2;
input 	temp_imemload_output_3;
input 	temp_imemload_output_5;
output 	Equal31;
input 	temp_imemload_output_15;
input 	temp_imemload_output_14;
input 	temp_imemload_output_13;
input 	temp_imemload_output_12;
input 	temp_imemload_output_11;
input 	temp_imemload_output_10;
input 	temp_imemload_output_9;
input 	temp_imemload_output_8;
input 	temp_imemload_output_7;
input 	temp_imemload_output_6;
input 	temp_imemload_output_1;
input 	temp_imemload_output_4;
output 	Equal32;
output 	WideOr8;
output 	WideOr2;
output 	WideOr4;
output 	WideOr7;
output 	WideOr1;
output 	WideOr5;
output 	WideOr6;
output 	WideOr0;
output 	halt_out;
output 	halt_out1;
output 	WideOr3;
output 	WideOr10;
output 	memtoreg;
output 	WideOr9;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Equal3~5_combout ;
wire \Equal3~6_combout ;
wire \Equal3~7_combout ;
wire \Equal3~4_combout ;
wire \Equal3~8_combout ;
wire \Equal3~2_combout ;
wire \Equal3~3_combout ;
wire \halt_out~1_combout ;
wire \halt_out~2_combout ;


// Location: LCCOMB_X65_Y40_N10
cycloneive_lcell_comb \Equal3~0 (
// Equation(s):
// Equal3 = (!temp_imemload_output_30 & (!temp_imemload_output_31 & (!temp_imemload_output_29 & !temp_imemload_output_28)))

	.dataa(temp_imemload_output_30),
	.datab(temp_imemload_output_31),
	.datac(temp_imemload_output_29),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(Equal3),
	.cout());
// synopsys translate_off
defparam \Equal3~0 .lut_mask = 16'h0001;
defparam \Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N6
cycloneive_lcell_comb \Equal3~1 (
// Equation(s):
// Equal31 = (!temp_imemload_output_0 & (!temp_imemload_output_5 & (!temp_imemload_output_2 & !temp_imemload_output_3)))

	.dataa(temp_imemload_output_0),
	.datab(temp_imemload_output_5),
	.datac(temp_imemload_output_2),
	.datad(temp_imemload_output_3),
	.cin(gnd),
	.combout(Equal31),
	.cout());
// synopsys translate_off
defparam \Equal3~1 .lut_mask = 16'h0001;
defparam \Equal3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N2
cycloneive_lcell_comb \Equal3~9 (
// Equation(s):
// Equal32 = (\Equal3~8_combout  & (!temp_imemload_output_1 & (!temp_imemload_output_4 & \Equal3~3_combout )))

	.dataa(\Equal3~8_combout ),
	.datab(temp_imemload_output_1),
	.datac(temp_imemload_output_4),
	.datad(\Equal3~3_combout ),
	.cin(gnd),
	.combout(Equal32),
	.cout());
// synopsys translate_off
defparam \Equal3~9 .lut_mask = 16'h0200;
defparam \Equal3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N4
cycloneive_lcell_comb \WideOr8~0 (
// Equation(s):
// WideOr8 = (temp_imemload_output_29 & (temp_imemload_output_26 & (temp_imemload_output_27 $ (temp_imemload_output_28)))) # (!temp_imemload_output_29 & (!temp_imemload_output_27 & ((temp_imemload_output_28))))

	.dataa(temp_imemload_output_27),
	.datab(temp_imemload_output_26),
	.datac(temp_imemload_output_29),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(WideOr8),
	.cout());
// synopsys translate_off
defparam \WideOr8~0 .lut_mask = 16'h4580;
defparam \WideOr8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N30
cycloneive_lcell_comb \WideOr2~0 (
// Equation(s):
// WideOr2 = (temp_imemload_output_0 & ((temp_imemload_output_2 & ((!temp_imemload_output_3))) # (!temp_imemload_output_2 & (temp_imemload_output_1))))

	.dataa(temp_imemload_output_0),
	.datab(temp_imemload_output_1),
	.datac(temp_imemload_output_2),
	.datad(temp_imemload_output_3),
	.cin(gnd),
	.combout(WideOr2),
	.cout());
// synopsys translate_off
defparam \WideOr2~0 .lut_mask = 16'h08A8;
defparam \WideOr2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N6
cycloneive_lcell_comb \WideOr4~0 (
// Equation(s):
// WideOr4 = (temp_imemload_output_27 & ((temp_imemload_output_26 & ((!temp_imemload_output_28))) # (!temp_imemload_output_26 & (!temp_imemload_output_31)))) # (!temp_imemload_output_27 & (!temp_imemload_output_31 & ((temp_imemload_output_26) # 
// (temp_imemload_output_28))))

	.dataa(temp_imemload_output_27),
	.datab(temp_imemload_output_31),
	.datac(temp_imemload_output_26),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(WideOr4),
	.cout());
// synopsys translate_off
defparam \WideOr4~0 .lut_mask = 16'h13B2;
defparam \WideOr4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N2
cycloneive_lcell_comb \WideOr7~0 (
// Equation(s):
// WideOr7 = (!temp_imemload_output_27 & ((temp_imemload_output_28) # ((temp_imemload_output_26 & temp_imemload_output_29))))

	.dataa(temp_imemload_output_27),
	.datab(temp_imemload_output_26),
	.datac(temp_imemload_output_29),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(WideOr7),
	.cout());
// synopsys translate_off
defparam \WideOr7~0 .lut_mask = 16'h5540;
defparam \WideOr7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N10
cycloneive_lcell_comb \WideOr1~0 (
// Equation(s):
// WideOr1 = (!temp_imemload_output_3 & ((temp_imemload_output_2 & ((!temp_imemload_output_1))) # (!temp_imemload_output_2 & (temp_imemload_output_0))))

	.dataa(temp_imemload_output_0),
	.datab(temp_imemload_output_1),
	.datac(temp_imemload_output_2),
	.datad(temp_imemload_output_3),
	.cin(gnd),
	.combout(WideOr1),
	.cout());
// synopsys translate_off
defparam \WideOr1~0 .lut_mask = 16'h003A;
defparam \WideOr1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N20
cycloneive_lcell_comb \WideOr5~0 (
// Equation(s):
// WideOr5 = (temp_imemload_output_29 & (!temp_imemload_output_28 & ((temp_imemload_output_27) # (temp_imemload_output_26)))) # (!temp_imemload_output_29 & (!temp_imemload_output_27 & ((temp_imemload_output_28))))

	.dataa(temp_imemload_output_27),
	.datab(temp_imemload_output_26),
	.datac(temp_imemload_output_29),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(WideOr5),
	.cout());
// synopsys translate_off
defparam \WideOr5~0 .lut_mask = 16'h05E0;
defparam \WideOr5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N14
cycloneive_lcell_comb \WideOr6~0 (
// Equation(s):
// WideOr6 = (temp_imemload_output_26 & (!temp_imemload_output_27 & (temp_imemload_output_29 $ (temp_imemload_output_28)))) # (!temp_imemload_output_26 & (temp_imemload_output_28 & (temp_imemload_output_27 $ (!temp_imemload_output_29))))

	.dataa(temp_imemload_output_27),
	.datab(temp_imemload_output_26),
	.datac(temp_imemload_output_29),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(WideOr6),
	.cout());
// synopsys translate_off
defparam \WideOr6~0 .lut_mask = 16'h2540;
defparam \WideOr6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N14
cycloneive_lcell_comb \WideOr0~0 (
// Equation(s):
// WideOr0 = (!temp_imemload_output_3 & ((temp_imemload_output_2 & ((temp_imemload_output_1))) # (!temp_imemload_output_2 & (temp_imemload_output_0))))

	.dataa(temp_imemload_output_0),
	.datab(temp_imemload_output_1),
	.datac(temp_imemload_output_2),
	.datad(temp_imemload_output_3),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
// synopsys translate_off
defparam \WideOr0~0 .lut_mask = 16'h00CA;
defparam \WideOr0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N28
cycloneive_lcell_comb \halt_out~0 (
// Equation(s):
// halt_out = (temp_imemload_output_3 & (temp_imemload_output_5 & temp_imemload_output_1))

	.dataa(gnd),
	.datab(temp_imemload_output_3),
	.datac(temp_imemload_output_5),
	.datad(temp_imemload_output_1),
	.cin(gnd),
	.combout(halt_out),
	.cout());
// synopsys translate_off
defparam \halt_out~0 .lut_mask = 16'hC000;
defparam \halt_out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N12
cycloneive_lcell_comb \halt_out~3 (
// Equation(s):
// halt_out1 = (\halt_out~1_combout  & (\halt_out~2_combout  & (temp_imemload_output_30 & halt_out)))

	.dataa(\halt_out~1_combout ),
	.datab(\halt_out~2_combout ),
	.datac(temp_imemload_output_30),
	.datad(halt_out),
	.cin(gnd),
	.combout(halt_out1),
	.cout());
// synopsys translate_off
defparam \halt_out~3 .lut_mask = 16'h8000;
defparam \halt_out~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N16
cycloneive_lcell_comb \WideOr3~0 (
// Equation(s):
// WideOr3 = (temp_imemload_output_2 & (((!temp_imemload_output_3)))) # (!temp_imemload_output_2 & ((temp_imemload_output_3 & ((temp_imemload_output_1))) # (!temp_imemload_output_3 & (temp_imemload_output_0))))

	.dataa(temp_imemload_output_0),
	.datab(temp_imemload_output_1),
	.datac(temp_imemload_output_2),
	.datad(temp_imemload_output_3),
	.cin(gnd),
	.combout(WideOr3),
	.cout());
// synopsys translate_off
defparam \WideOr3~0 .lut_mask = 16'h0CFA;
defparam \WideOr3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N24
cycloneive_lcell_comb \WideOr10~0 (
// Equation(s):
// WideOr10 = (temp_imemload_output_27 & ((temp_imemload_output_29) # ((temp_imemload_output_26 & !temp_imemload_output_28)))) # (!temp_imemload_output_27 & (temp_imemload_output_29 & ((temp_imemload_output_26) # (temp_imemload_output_28))))

	.dataa(temp_imemload_output_27),
	.datab(temp_imemload_output_26),
	.datac(temp_imemload_output_29),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(WideOr10),
	.cout());
// synopsys translate_off
defparam \WideOr10~0 .lut_mask = 16'hF0E8;
defparam \WideOr10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N2
cycloneive_lcell_comb \memtoreg~0 (
// Equation(s):
// memtoreg = (temp_imemload_output_27 & (temp_imemload_output_26 & (temp_imemload_output_29 $ (!temp_imemload_output_28))))

	.dataa(temp_imemload_output_27),
	.datab(temp_imemload_output_26),
	.datac(temp_imemload_output_29),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(memtoreg),
	.cout());
// synopsys translate_off
defparam \memtoreg~0 .lut_mask = 16'h8008;
defparam \memtoreg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N22
cycloneive_lcell_comb \WideOr9~0 (
// Equation(s):
// WideOr9 = (!temp_imemload_output_29 & (!temp_imemload_output_30 & (temp_imemload_output_27 $ (temp_imemload_output_28))))

	.dataa(temp_imemload_output_27),
	.datab(temp_imemload_output_29),
	.datac(temp_imemload_output_30),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(WideOr9),
	.cout());
// synopsys translate_off
defparam \WideOr9~0 .lut_mask = 16'h0102;
defparam \WideOr9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N16
cycloneive_lcell_comb \Equal3~5 (
// Equation(s):
// \Equal3~5_combout  = (!temp_imemload_output_14 & (!temp_imemload_output_15 & (!temp_imemload_output_17 & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_14),
	.datab(temp_imemload_output_15),
	.datac(temp_imemload_output_17),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Equal3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~5 .lut_mask = 16'h0001;
defparam \Equal3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N14
cycloneive_lcell_comb \Equal3~6 (
// Equation(s):
// \Equal3~6_combout  = (!temp_imemload_output_13 & (!temp_imemload_output_12 & (!temp_imemload_output_11 & !temp_imemload_output_10)))

	.dataa(temp_imemload_output_13),
	.datab(temp_imemload_output_12),
	.datac(temp_imemload_output_11),
	.datad(temp_imemload_output_10),
	.cin(gnd),
	.combout(\Equal3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~6 .lut_mask = 16'h0001;
defparam \Equal3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N24
cycloneive_lcell_comb \Equal3~7 (
// Equation(s):
// \Equal3~7_combout  = (!temp_imemload_output_8 & (!temp_imemload_output_9 & (!temp_imemload_output_6 & !temp_imemload_output_7)))

	.dataa(temp_imemload_output_8),
	.datab(temp_imemload_output_9),
	.datac(temp_imemload_output_6),
	.datad(temp_imemload_output_7),
	.cin(gnd),
	.combout(\Equal3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~7 .lut_mask = 16'h0001;
defparam \Equal3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N24
cycloneive_lcell_comb \Equal3~4 (
// Equation(s):
// \Equal3~4_combout  = (!temp_imemload_output_21 & (!temp_imemload_output_18 & (!temp_imemload_output_20 & !temp_imemload_output_19)))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_18),
	.datac(temp_imemload_output_20),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Equal3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~4 .lut_mask = 16'h0001;
defparam \Equal3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N10
cycloneive_lcell_comb \Equal3~8 (
// Equation(s):
// \Equal3~8_combout  = (\Equal3~5_combout  & (\Equal3~6_combout  & (\Equal3~7_combout  & \Equal3~4_combout )))

	.dataa(\Equal3~5_combout ),
	.datab(\Equal3~6_combout ),
	.datac(\Equal3~7_combout ),
	.datad(\Equal3~4_combout ),
	.cin(gnd),
	.combout(\Equal3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~8 .lut_mask = 16'h8000;
defparam \Equal3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N0
cycloneive_lcell_comb \Equal3~2 (
// Equation(s):
// \Equal3~2_combout  = (!temp_imemload_output_25 & (!temp_imemload_output_22 & (!temp_imemload_output_23 & !temp_imemload_output_24)))

	.dataa(temp_imemload_output_25),
	.datab(temp_imemload_output_22),
	.datac(temp_imemload_output_23),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Equal3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~2 .lut_mask = 16'h0001;
defparam \Equal3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N0
cycloneive_lcell_comb \Equal3~3 (
// Equation(s):
// \Equal3~3_combout  = (Equal31 & (Equal3 & (temp_branch_output1 & \Equal3~2_combout )))

	.dataa(Equal31),
	.datab(Equal3),
	.datac(temp_branch_output),
	.datad(\Equal3~2_combout ),
	.cin(gnd),
	.combout(\Equal3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~3 .lut_mask = 16'h8000;
defparam \Equal3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N10
cycloneive_lcell_comb \halt_out~1 (
// Equation(s):
// \halt_out~1_combout  = (temp_imemload_output_27 & (temp_imemload_output_0 & (temp_imemload_output_26 & temp_imemload_output_31)))

	.dataa(temp_imemload_output_27),
	.datab(temp_imemload_output_0),
	.datac(temp_imemload_output_26),
	.datad(temp_imemload_output_31),
	.cin(gnd),
	.combout(\halt_out~1_combout ),
	.cout());
// synopsys translate_off
defparam \halt_out~1 .lut_mask = 16'h8000;
defparam \halt_out~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N20
cycloneive_lcell_comb \halt_out~2 (
// Equation(s):
// \halt_out~2_combout  = (temp_imemload_output_4 & (temp_imemload_output_29 & (temp_imemload_output_2 & temp_imemload_output_28)))

	.dataa(temp_imemload_output_4),
	.datab(temp_imemload_output_29),
	.datac(temp_imemload_output_2),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(\halt_out~2_combout ),
	.cout());
// synopsys translate_off
defparam \halt_out~2 .lut_mask = 16'h8000;
defparam \halt_out~2 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module ex_mem_latch (
	temp_branchDest_0,
	temp_branchDest_4,
	temp_branchDest_3,
	temp_branchDest_2,
	temp_branchDest_1,
	temp_signzerovalue_output_16,
	temp_zeroFlag1,
	temp_halt_out_output,
	temp_aluResult_1,
	temp_dmemWEN1,
	temp_dmemREN1,
	temp_aluResult_0,
	temp_aluResult_2,
	temp_aluResult_3,
	temp_aluResult_5,
	temp_aluResult_4,
	temp_aluResult_7,
	temp_aluResult_6,
	temp_aluResult_9,
	temp_aluResult_8,
	temp_aluResult_11,
	temp_aluResult_10,
	temp_aluResult_13,
	temp_aluResult_12,
	temp_aluResult_15,
	temp_aluResult_14,
	temp_aluResult_17,
	temp_aluResult_16,
	temp_aluResult_19,
	temp_aluResult_18,
	temp_aluResult_20,
	temp_aluResult_21,
	temp_aluResult_23,
	temp_aluResult_22,
	temp_aluResult_25,
	temp_aluResult_24,
	temp_aluResult_26,
	temp_aluResult_27,
	temp_aluResult_29,
	temp_aluResult_28,
	temp_aluResult_31,
	temp_aluResult_30,
	temp_halt_out1,
	temp_rdat2_0,
	temp_imemload_output_1,
	temp_imemload_output_7,
	temp_regwrite1,
	temp_imemload_output_17,
	temp_imemload_output_16,
	temp_imemload_output_18,
	temp_imemload_output_19,
	temp_imemload_output_20,
	temp_memtoreg_0,
	temp_memtoreg_1,
	alu_b_mux_output_1,
	alu_b_mux_output_11,
	temp_imemload_output_22,
	temp_imemload_output_21,
	temp_imemload_output_23,
	alu_a_mux_output_1,
	alu_b_mux_output_0,
	temp_imemload_output_0,
	temp_imemload_output_6,
	alu_b_mux_output_01,
	alu_a_mux_output_0,
	alu_a_mux_output_2,
	alu_a_mux_output_4,
	alu_a_mux_output_3,
	temp_imemload_output_2,
	temp_imemload_output_8,
	alu_b_mux_output_2,
	alu_a_mux_output_8,
	alu_a_mux_output_7,
	alu_a_mux_output_6,
	alu_a_mux_output_5,
	temp_imemload_output_3,
	temp_imemload_output_9,
	alu_b_mux_output_3,
	temp_iMemLoad_0,
	alu_a_mux_output_16,
	alu_a_mux_output_14,
	alu_a_mux_output_15,
	alu_a_mux_output_13,
	alu_a_mux_output_12,
	alu_a_mux_output_10,
	alu_a_mux_output_11,
	alu_a_mux_output_9,
	temp_imemload_output_4,
	temp_imemload_output_10,
	alu_b_mux_output_4,
	temp_iMemLoad_15,
	alu_a_mux_output_31,
	temp_iMemLoad_14,
	alu_a_mux_output_30,
	temp_iMemLoad_13,
	alu_a_mux_output_29,
	temp_iMemLoad_10,
	alu_a_mux_output_26,
	temp_iMemLoad_9,
	alu_a_mux_output_25,
	temp_iMemLoad_12,
	alu_a_mux_output_28,
	temp_iMemLoad_11,
	alu_a_mux_output_27,
	temp_iMemLoad_1,
	alu_a_mux_output_17,
	temp_iMemLoad_4,
	alu_a_mux_output_20,
	temp_iMemLoad_3,
	alu_a_mux_output_19,
	temp_iMemLoad_2,
	alu_a_mux_output_18,
	temp_iMemLoad_8,
	alu_a_mux_output_24,
	temp_iMemLoad_7,
	alu_a_mux_output_23,
	temp_iMemLoad_6,
	alu_a_mux_output_22,
	temp_iMemLoad_5,
	alu_a_mux_output_21,
	alu_b_mux_output_15,
	temp_imemload_output_15,
	alu_b_mux_output_12,
	temp_imemload_output_12,
	alu_b_mux_output_27,
	alu_b_mux_output_18,
	alu_b_mux_output_17,
	alu_b_mux_output_16,
	alu_b_mux_output_31,
	alu_b_mux_output_30,
	alu_b_mux_output_29,
	alu_b_mux_output_28,
	alu_b_mux_output_26,
	alu_b_mux_output_25,
	alu_b_mux_output_24,
	alu_b_mux_output_23,
	alu_b_mux_output_22,
	alu_b_mux_output_21,
	alu_b_mux_output_20,
	alu_b_mux_output_19,
	temp_imemload_output_14,
	alu_b_mux_output_10,
	alu_b_mux_output_14,
	alu_b_mux_output_9,
	alu_b_mux_output_8,
	alu_b_mux_output_7,
	alu_b_mux_output_6,
	alu_b_mux_output_5,
	temp_imemload_output_5,
	alu_b_mux_output_13,
	temp_imemload_output_13,
	alu_b_mux_output_111,
	temp_imemload_output_11,
	temp_ALUop_output_3,
	Mux30,
	temp_iMemLoad_31,
	temp_iMemLoad_30,
	temp_iMemLoad_29,
	ex_mem_flush,
	temp_iMemLoad_27,
	temp_iMemLoad_26,
	temp_iMemLoad_28,
	ex_mem_flush1,
	temp_branchSelect1,
	ex_mem_flush2,
	ex_mem_flush3,
	wen,
	temp_rdat1_1,
	temp_npc_1,
	temp_pcselect_1,
	temp_pcselect_0,
	temp_request_dmemREN_output,
	temp_request_dmemWEN_output,
	Mux31,
	temp_rdat1_0,
	temp_npc_0,
	Mux29,
	temp_npc_2,
	temp_rdat1_2,
	Mux28,
	temp_npc_3,
	temp_rdat1_3,
	alu_a_mux_output_32,
	Mux26,
	temp_npc_5,
	temp_npc_4,
	temp_rdat1_5,
	Mux27,
	temp_rdat1_4,
	Mux24,
	temp_npc_7,
	temp_npc_6,
	temp_rdat1_7,
	Mux25,
	temp_rdat1_6,
	Mux22,
	Mux221,
	Mux19,
	temp_npc_9,
	temp_npc_8,
	temp_rdat1_9,
	Mux23,
	Mux231,
	temp_rdat1_8,
	Mux20,
	Mux201,
	temp_npc_11,
	temp_npc_10,
	temp_rdat1_11,
	Mux21,
	Mux211,
	temp_rdat1_10,
	Mux18,
	Mux181,
	temp_npc_13,
	temp_npc_12,
	temp_rdat1_13,
	Mux191,
	Mux192,
	temp_rdat1_12,
	Mux16,
	Mux161,
	temp_npc_15,
	temp_npc_14,
	temp_rdat1_15,
	Mux17,
	Mux171,
	temp_rdat1_14,
	Mux14,
	Mux141,
	temp_npc_17,
	temp_npc_16,
	temp_rdat1_17,
	Mux15,
	Mux151,
	temp_rdat1_16,
	Mux12,
	Mux121,
	temp_signZero_16,
	temp_npc_19,
	temp_npc_18,
	temp_rdat1_19,
	temp_iMemLoad_17,
	Mux13,
	Mux131,
	temp_rdat1_18,
	temp_iMemLoad_16,
	Mux11,
	Mux111,
	temp_npc_20,
	temp_rdat1_20,
	temp_iMemLoad_18,
	Mux10,
	Mux101,
	temp_npc_21,
	temp_rdat1_21,
	temp_iMemLoad_19,
	Mux8,
	Mux81,
	temp_npc_23,
	temp_npc_22,
	temp_rdat1_23,
	temp_iMemLoad_21,
	Mux9,
	Mux91,
	temp_rdat1_22,
	temp_iMemLoad_20,
	Mux6,
	temp_npc_25,
	temp_npc_24,
	temp_rdat1_25,
	temp_iMemLoad_23,
	temp_rdat1_24,
	temp_iMemLoad_22,
	temp_npc_26,
	temp_rdat1_26,
	Mux4,
	temp_npc_27,
	temp_rdat1_27,
	Mux2,
	temp_npc_29,
	temp_npc_28,
	temp_rdat1_29,
	Mux3,
	temp_rdat1_28,
	Mux0,
	Mux01,
	temp_rdat1_31,
	temp_npc_31,
	temp_npc_30,
	Mux1,
	temp_rdat1_30,
	temp_rdat2_1,
	temp_rdat2_2,
	temp_rdat2_3,
	temp_rdat2_4,
	temp_rdat2_5,
	temp_rdat2_6,
	temp_rdat2_7,
	temp_rdat2_8,
	temp_rdat2_9,
	temp_rdat2_10,
	temp_rdat2_11,
	temp_rdat2_12,
	temp_rdat2_13,
	temp_rdat2_14,
	temp_rdat2_15,
	temp_rdat2_16,
	temp_rdat2_17,
	temp_rdat2_18,
	temp_rdat2_19,
	temp_rdat2_20,
	temp_rdat2_21,
	temp_rdat2_22,
	temp_rdat2_23,
	temp_rdat2_24,
	temp_rdat2_25,
	temp_rdat2_26,
	temp_rdat2_27,
	temp_rdat2_28,
	temp_rdat2_29,
	temp_rdat2_30,
	temp_rdat2_31,
	temp_regwrite_output,
	temp_regdst_output_1,
	temp_regdst_output_0,
	temp_memtoreg_output_0,
	temp_memtoreg_output_1,
	temp_imemload_output_31,
	temp_imemload_output_30,
	temp_imemload_output_29,
	temp_imemload_output_27,
	temp_imemload_output_26,
	temp_imemload_output_28,
	temp_branch_output,
	Equal0,
	temp_NPC_output_1,
	temp_pcselect_output_1,
	temp_pcselect_output_0,
	temp_NPC_output_0,
	temp_NPC_output_2,
	temp_NPC_output_3,
	temp_NPC_output_5,
	temp_NPC_output_4,
	temp_NPC_output_7,
	temp_NPC_output_6,
	temp_NPC_output_9,
	temp_NPC_output_8,
	temp_NPC_output_11,
	temp_NPC_output_10,
	temp_NPC_output_13,
	temp_NPC_output_12,
	temp_NPC_output_15,
	temp_NPC_output_14,
	temp_NPC_output_17,
	temp_NPC_output_16,
	temp_NPC_output_19,
	temp_NPC_output_18,
	temp_NPC_output_20,
	temp_NPC_output_21,
	temp_NPC_output_23,
	temp_NPC_output_22,
	temp_NPC_output_25,
	temp_NPC_output_24,
	temp_NPC_output_26,
	temp_NPC_output_27,
	temp_NPC_output_29,
	temp_NPC_output_28,
	temp_NPC_output_31,
	temp_NPC_output_30,
	Mux110,
	Mux5,
	Mux7,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	temp_branchDest_0;
output 	temp_branchDest_4;
output 	temp_branchDest_3;
output 	temp_branchDest_2;
output 	temp_branchDest_1;
input 	temp_signzerovalue_output_16;
output 	temp_zeroFlag1;
input 	temp_halt_out_output;
output 	temp_aluResult_1;
output 	temp_dmemWEN1;
output 	temp_dmemREN1;
output 	temp_aluResult_0;
output 	temp_aluResult_2;
output 	temp_aluResult_3;
output 	temp_aluResult_5;
output 	temp_aluResult_4;
output 	temp_aluResult_7;
output 	temp_aluResult_6;
output 	temp_aluResult_9;
output 	temp_aluResult_8;
output 	temp_aluResult_11;
output 	temp_aluResult_10;
output 	temp_aluResult_13;
output 	temp_aluResult_12;
output 	temp_aluResult_15;
output 	temp_aluResult_14;
output 	temp_aluResult_17;
output 	temp_aluResult_16;
output 	temp_aluResult_19;
output 	temp_aluResult_18;
output 	temp_aluResult_20;
output 	temp_aluResult_21;
output 	temp_aluResult_23;
output 	temp_aluResult_22;
output 	temp_aluResult_25;
output 	temp_aluResult_24;
output 	temp_aluResult_26;
output 	temp_aluResult_27;
output 	temp_aluResult_29;
output 	temp_aluResult_28;
output 	temp_aluResult_31;
output 	temp_aluResult_30;
output 	temp_halt_out1;
output 	temp_rdat2_0;
input 	temp_imemload_output_1;
input 	temp_imemload_output_7;
output 	temp_regwrite1;
input 	temp_imemload_output_17;
input 	temp_imemload_output_16;
input 	temp_imemload_output_18;
input 	temp_imemload_output_19;
input 	temp_imemload_output_20;
output 	temp_memtoreg_0;
output 	temp_memtoreg_1;
input 	alu_b_mux_output_1;
input 	alu_b_mux_output_11;
input 	temp_imemload_output_22;
input 	temp_imemload_output_21;
input 	temp_imemload_output_23;
input 	alu_a_mux_output_1;
input 	alu_b_mux_output_0;
input 	temp_imemload_output_0;
input 	temp_imemload_output_6;
input 	alu_b_mux_output_01;
input 	alu_a_mux_output_0;
input 	alu_a_mux_output_2;
input 	alu_a_mux_output_4;
input 	alu_a_mux_output_3;
input 	temp_imemload_output_2;
input 	temp_imemload_output_8;
input 	alu_b_mux_output_2;
input 	alu_a_mux_output_8;
input 	alu_a_mux_output_7;
input 	alu_a_mux_output_6;
input 	alu_a_mux_output_5;
input 	temp_imemload_output_3;
input 	temp_imemload_output_9;
input 	alu_b_mux_output_3;
output 	temp_iMemLoad_0;
input 	alu_a_mux_output_16;
input 	alu_a_mux_output_14;
input 	alu_a_mux_output_15;
input 	alu_a_mux_output_13;
input 	alu_a_mux_output_12;
input 	alu_a_mux_output_10;
input 	alu_a_mux_output_11;
input 	alu_a_mux_output_9;
input 	temp_imemload_output_4;
input 	temp_imemload_output_10;
input 	alu_b_mux_output_4;
output 	temp_iMemLoad_15;
input 	alu_a_mux_output_31;
output 	temp_iMemLoad_14;
input 	alu_a_mux_output_30;
output 	temp_iMemLoad_13;
input 	alu_a_mux_output_29;
output 	temp_iMemLoad_10;
input 	alu_a_mux_output_26;
output 	temp_iMemLoad_9;
input 	alu_a_mux_output_25;
output 	temp_iMemLoad_12;
input 	alu_a_mux_output_28;
output 	temp_iMemLoad_11;
input 	alu_a_mux_output_27;
output 	temp_iMemLoad_1;
input 	alu_a_mux_output_17;
output 	temp_iMemLoad_4;
input 	alu_a_mux_output_20;
output 	temp_iMemLoad_3;
input 	alu_a_mux_output_19;
output 	temp_iMemLoad_2;
input 	alu_a_mux_output_18;
output 	temp_iMemLoad_8;
input 	alu_a_mux_output_24;
output 	temp_iMemLoad_7;
input 	alu_a_mux_output_23;
output 	temp_iMemLoad_6;
input 	alu_a_mux_output_22;
output 	temp_iMemLoad_5;
input 	alu_a_mux_output_21;
input 	alu_b_mux_output_15;
input 	temp_imemload_output_15;
input 	alu_b_mux_output_12;
input 	temp_imemload_output_12;
input 	alu_b_mux_output_27;
input 	alu_b_mux_output_18;
input 	alu_b_mux_output_17;
input 	alu_b_mux_output_16;
input 	alu_b_mux_output_31;
input 	alu_b_mux_output_30;
input 	alu_b_mux_output_29;
input 	alu_b_mux_output_28;
input 	alu_b_mux_output_26;
input 	alu_b_mux_output_25;
input 	alu_b_mux_output_24;
input 	alu_b_mux_output_23;
input 	alu_b_mux_output_22;
input 	alu_b_mux_output_21;
input 	alu_b_mux_output_20;
input 	alu_b_mux_output_19;
input 	temp_imemload_output_14;
input 	alu_b_mux_output_10;
input 	alu_b_mux_output_14;
input 	alu_b_mux_output_9;
input 	alu_b_mux_output_8;
input 	alu_b_mux_output_7;
input 	alu_b_mux_output_6;
input 	alu_b_mux_output_5;
input 	temp_imemload_output_5;
input 	alu_b_mux_output_13;
input 	temp_imemload_output_13;
input 	alu_b_mux_output_111;
input 	temp_imemload_output_11;
input 	temp_ALUop_output_3;
input 	Mux30;
output 	temp_iMemLoad_31;
output 	temp_iMemLoad_30;
output 	temp_iMemLoad_29;
input 	ex_mem_flush;
output 	temp_iMemLoad_27;
output 	temp_iMemLoad_26;
output 	temp_iMemLoad_28;
input 	ex_mem_flush1;
output 	temp_branchSelect1;
input 	ex_mem_flush2;
input 	ex_mem_flush3;
input 	wen;
output 	temp_rdat1_1;
output 	temp_npc_1;
output 	temp_pcselect_1;
output 	temp_pcselect_0;
input 	temp_request_dmemREN_output;
input 	temp_request_dmemWEN_output;
input 	Mux31;
output 	temp_rdat1_0;
output 	temp_npc_0;
input 	Mux29;
output 	temp_npc_2;
output 	temp_rdat1_2;
input 	Mux28;
output 	temp_npc_3;
output 	temp_rdat1_3;
input 	alu_a_mux_output_32;
input 	Mux26;
output 	temp_npc_5;
output 	temp_npc_4;
output 	temp_rdat1_5;
input 	Mux27;
output 	temp_rdat1_4;
input 	Mux24;
output 	temp_npc_7;
output 	temp_npc_6;
output 	temp_rdat1_7;
input 	Mux25;
output 	temp_rdat1_6;
input 	Mux22;
input 	Mux221;
input 	Mux19;
output 	temp_npc_9;
output 	temp_npc_8;
output 	temp_rdat1_9;
input 	Mux23;
input 	Mux231;
output 	temp_rdat1_8;
input 	Mux20;
input 	Mux201;
output 	temp_npc_11;
output 	temp_npc_10;
output 	temp_rdat1_11;
input 	Mux21;
input 	Mux211;
output 	temp_rdat1_10;
input 	Mux18;
input 	Mux181;
output 	temp_npc_13;
output 	temp_npc_12;
output 	temp_rdat1_13;
input 	Mux191;
input 	Mux192;
output 	temp_rdat1_12;
input 	Mux16;
input 	Mux161;
output 	temp_npc_15;
output 	temp_npc_14;
output 	temp_rdat1_15;
input 	Mux17;
input 	Mux171;
output 	temp_rdat1_14;
input 	Mux14;
input 	Mux141;
output 	temp_npc_17;
output 	temp_npc_16;
output 	temp_rdat1_17;
input 	Mux15;
input 	Mux151;
output 	temp_rdat1_16;
input 	Mux12;
input 	Mux121;
output 	temp_signZero_16;
output 	temp_npc_19;
output 	temp_npc_18;
output 	temp_rdat1_19;
output 	temp_iMemLoad_17;
input 	Mux13;
input 	Mux131;
output 	temp_rdat1_18;
output 	temp_iMemLoad_16;
input 	Mux11;
input 	Mux111;
output 	temp_npc_20;
output 	temp_rdat1_20;
output 	temp_iMemLoad_18;
input 	Mux10;
input 	Mux101;
output 	temp_npc_21;
output 	temp_rdat1_21;
output 	temp_iMemLoad_19;
input 	Mux8;
input 	Mux81;
output 	temp_npc_23;
output 	temp_npc_22;
output 	temp_rdat1_23;
output 	temp_iMemLoad_21;
input 	Mux9;
input 	Mux91;
output 	temp_rdat1_22;
output 	temp_iMemLoad_20;
input 	Mux6;
output 	temp_npc_25;
output 	temp_npc_24;
output 	temp_rdat1_25;
output 	temp_iMemLoad_23;
output 	temp_rdat1_24;
output 	temp_iMemLoad_22;
output 	temp_npc_26;
output 	temp_rdat1_26;
input 	Mux4;
output 	temp_npc_27;
output 	temp_rdat1_27;
input 	Mux2;
output 	temp_npc_29;
output 	temp_npc_28;
output 	temp_rdat1_29;
input 	Mux3;
output 	temp_rdat1_28;
input 	Mux0;
input 	Mux01;
output 	temp_rdat1_31;
output 	temp_npc_31;
output 	temp_npc_30;
input 	Mux1;
output 	temp_rdat1_30;
output 	temp_rdat2_1;
output 	temp_rdat2_2;
output 	temp_rdat2_3;
output 	temp_rdat2_4;
output 	temp_rdat2_5;
output 	temp_rdat2_6;
output 	temp_rdat2_7;
output 	temp_rdat2_8;
output 	temp_rdat2_9;
output 	temp_rdat2_10;
output 	temp_rdat2_11;
output 	temp_rdat2_12;
output 	temp_rdat2_13;
output 	temp_rdat2_14;
output 	temp_rdat2_15;
output 	temp_rdat2_16;
output 	temp_rdat2_17;
output 	temp_rdat2_18;
output 	temp_rdat2_19;
output 	temp_rdat2_20;
output 	temp_rdat2_21;
output 	temp_rdat2_22;
output 	temp_rdat2_23;
output 	temp_rdat2_24;
output 	temp_rdat2_25;
output 	temp_rdat2_26;
output 	temp_rdat2_27;
output 	temp_rdat2_28;
output 	temp_rdat2_29;
output 	temp_rdat2_30;
output 	temp_rdat2_31;
input 	temp_regwrite_output;
input 	temp_regdst_output_1;
input 	temp_regdst_output_0;
input 	temp_memtoreg_output_0;
input 	temp_memtoreg_output_1;
input 	temp_imemload_output_31;
input 	temp_imemload_output_30;
input 	temp_imemload_output_29;
input 	temp_imemload_output_27;
input 	temp_imemload_output_26;
input 	temp_imemload_output_28;
input 	temp_branch_output;
input 	Equal0;
input 	temp_NPC_output_1;
input 	temp_pcselect_output_1;
input 	temp_pcselect_output_0;
input 	temp_NPC_output_0;
input 	temp_NPC_output_2;
input 	temp_NPC_output_3;
input 	temp_NPC_output_5;
input 	temp_NPC_output_4;
input 	temp_NPC_output_7;
input 	temp_NPC_output_6;
input 	temp_NPC_output_9;
input 	temp_NPC_output_8;
input 	temp_NPC_output_11;
input 	temp_NPC_output_10;
input 	temp_NPC_output_13;
input 	temp_NPC_output_12;
input 	temp_NPC_output_15;
input 	temp_NPC_output_14;
input 	temp_NPC_output_17;
input 	temp_NPC_output_16;
input 	temp_NPC_output_19;
input 	temp_NPC_output_18;
input 	temp_NPC_output_20;
input 	temp_NPC_output_21;
input 	temp_NPC_output_23;
input 	temp_NPC_output_22;
input 	temp_NPC_output_25;
input 	temp_NPC_output_24;
input 	temp_NPC_output_26;
input 	temp_NPC_output_27;
input 	temp_NPC_output_29;
input 	temp_NPC_output_28;
input 	temp_NPC_output_31;
input 	temp_NPC_output_30;
input 	Mux110;
input 	Mux5;
input 	Mux7;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \temp_branchDest~0_combout ;
wire \temp_branchDest~1_combout ;
wire \temp_branchDest~2_combout ;
wire \temp_branchDest~3_combout ;
wire \temp_branchDest~4_combout ;
wire \temp_aluResult~35_combout ;
wire \temp_dmemWEN~0_combout ;
wire \temp_dmemWEN~feeder_combout ;
wire \temp_dmemREN~0_combout ;
wire \temp_dmemREN~feeder_combout ;
wire \temp_aluResult~36_combout ;
wire \temp_aluResult~4_combout ;
wire \temp_aluResult~5_combout ;
wire \temp_aluResult~6_combout ;
wire \temp_aluResult~7_combout ;
wire \temp_aluResult~8_combout ;
wire \temp_aluResult~9_combout ;
wire \temp_aluResult~10_combout ;
wire \temp_aluResult~11_combout ;
wire \temp_aluResult~12_combout ;
wire \temp_aluResult~13_combout ;
wire \temp_aluResult~14_combout ;
wire \temp_aluResult~15_combout ;
wire \temp_aluResult~16_combout ;
wire \temp_aluResult~17_combout ;
wire \temp_aluResult~18_combout ;
wire \temp_aluResult~19_combout ;
wire \temp_aluResult~20_combout ;
wire \temp_aluResult~21_combout ;
wire \temp_aluResult~22_combout ;
wire \temp_aluResult~23_combout ;
wire \temp_aluResult~24_combout ;
wire \temp_aluResult~25_combout ;
wire \temp_aluResult~26_combout ;
wire \temp_aluResult~27_combout ;
wire \temp_aluResult~28_combout ;
wire \temp_aluResult~29_combout ;
wire \temp_aluResult~30_combout ;
wire \temp_aluResult~31_combout ;
wire \temp_aluResult~32_combout ;
wire \temp_aluResult~33_combout ;
wire \temp_aluResult~34_combout ;
wire \temp_halt_out~0_combout ;
wire \temp_rdat2~60_combout ;
wire \temp_regwrite~0_combout ;
wire \temp_memtoreg~0_combout ;
wire \temp_memtoreg~1_combout ;
wire \temp_iMemLoad~0_combout ;
wire \temp_iMemLoad~1_combout ;
wire \temp_iMemLoad~2_combout ;
wire \temp_iMemLoad~3_combout ;
wire \temp_iMemLoad~4_combout ;
wire \temp_iMemLoad~5_combout ;
wire \temp_iMemLoad~6_combout ;
wire \temp_iMemLoad~7_combout ;
wire \temp_iMemLoad~8_combout ;
wire \temp_iMemLoad~9_combout ;
wire \temp_iMemLoad~10_combout ;
wire \temp_iMemLoad~11_combout ;
wire \temp_iMemLoad~12_combout ;
wire \temp_iMemLoad~13_combout ;
wire \temp_iMemLoad~14_combout ;
wire \temp_iMemLoad~15_combout ;
wire \temp_iMemLoad~16_combout ;
wire \temp_iMemLoad~17_combout ;
wire \temp_iMemLoad~18_combout ;
wire \temp_iMemLoad~19_combout ;
wire \temp_iMemLoad~20_combout ;
wire \temp_iMemLoad~21_combout ;
wire \temp_branchSelect~0_combout ;
wire \temp_rdat1~63_combout ;
wire \temp_npc~0_combout ;
wire \temp_pcselect~0_combout ;
wire \temp_pcselect~1_combout ;
wire \temp_rdat1~64_combout ;
wire \temp_npc~1_combout ;
wire \temp_npc~2_combout ;
wire \temp_rdat1~65_combout ;
wire \temp_npc~3_combout ;
wire \temp_rdat1~62_combout ;
wire \temp_npc~4_combout ;
wire \temp_npc~5_combout ;
wire \temp_rdat1~66_combout ;
wire \temp_rdat1~67_combout ;
wire \temp_npc~6_combout ;
wire \temp_npc~7_combout ;
wire \temp_rdat1~68_combout ;
wire \temp_rdat1~69_combout ;
wire \temp_rdat1[6]~feeder_combout ;
wire \temp_npc~8_combout ;
wire \temp_npc~9_combout ;
wire \temp_rdat1~70_combout ;
wire \temp_rdat1~71_combout ;
wire \temp_npc~10_combout ;
wire \temp_npc~11_combout ;
wire \temp_rdat1~72_combout ;
wire \temp_rdat1~73_combout ;
wire \temp_npc~12_combout ;
wire \temp_npc~13_combout ;
wire \temp_rdat1~74_combout ;
wire \temp_rdat1~75_combout ;
wire \temp_npc~14_combout ;
wire \temp_npc~15_combout ;
wire \temp_rdat1~76_combout ;
wire \temp_rdat1~77_combout ;
wire \temp_npc~16_combout ;
wire \temp_npc~17_combout ;
wire \temp_rdat1~78_combout ;
wire \temp_rdat1~79_combout ;
wire \temp_signZero~0_combout ;
wire \temp_npc~18_combout ;
wire \temp_npc~19_combout ;
wire \temp_rdat1~80_combout ;
wire \temp_iMemLoad~22_combout ;
wire \temp_rdat1~81_combout ;
wire \temp_iMemLoad~23_combout ;
wire \temp_npc~20_combout ;
wire \temp_rdat1~82_combout ;
wire \temp_iMemLoad~24_combout ;
wire \temp_npc~21_combout ;
wire \temp_rdat1~83_combout ;
wire \temp_iMemLoad~25_combout ;
wire \temp_npc~22_combout ;
wire \temp_npc~23_combout ;
wire \temp_rdat1~84_combout ;
wire \temp_iMemLoad~26_combout ;
wire \temp_rdat1~85_combout ;
wire \temp_iMemLoad~27_combout ;
wire \temp_npc~24_combout ;
wire \temp_npc~25_combout ;
wire \temp_rdat1~86_combout ;
wire \temp_iMemLoad~28_combout ;
wire \temp_rdat1~87_combout ;
wire \temp_iMemLoad~29_combout ;
wire \temp_npc~26_combout ;
wire \temp_rdat1~88_combout ;
wire \temp_npc~27_combout ;
wire \temp_rdat1~89_combout ;
wire \temp_npc~28_combout ;
wire \temp_npc~29_combout ;
wire \temp_rdat1~90_combout ;
wire \temp_rdat1~91_combout ;
wire \temp_rdat1~92_combout ;
wire \temp_npc~30_combout ;
wire \temp_npc~31_combout ;
wire \temp_rdat1~93_combout ;
wire \temp_rdat2~61_combout ;
wire \temp_rdat2~62_combout ;
wire \temp_rdat2~63_combout ;
wire \temp_rdat2~64_combout ;
wire \temp_rdat2~65_combout ;
wire \temp_rdat2~66_combout ;
wire \temp_rdat2~67_combout ;
wire \temp_rdat2~68_combout ;
wire \temp_rdat2~69_combout ;
wire \temp_rdat2~70_combout ;
wire \temp_rdat2~71_combout ;
wire \temp_rdat2~72_combout ;
wire \temp_rdat2~73_combout ;
wire \temp_rdat2~74_combout ;
wire \temp_rdat2~75_combout ;
wire \temp_rdat2~76_combout ;
wire \temp_rdat2~77_combout ;
wire \temp_rdat2~78_combout ;
wire \temp_rdat2~79_combout ;
wire \temp_rdat2~80_combout ;
wire \temp_rdat2~81_combout ;
wire \temp_rdat2~82_combout ;
wire \temp_rdat2~83_combout ;
wire \temp_rdat2~84_combout ;
wire \temp_rdat2~85_combout ;
wire \temp_rdat2~86_combout ;
wire \temp_rdat2~87_combout ;
wire \temp_rdat2~88_combout ;
wire \temp_rdat2~89_combout ;
wire \temp_rdat2~90_combout ;
wire \temp_rdat2~91_combout ;


// Location: FF_X59_Y41_N5
dffeas \temp_branchDest[0] (
	.clk(CLK),
	.d(\temp_branchDest~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(ex_mem_flush3),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branchDest_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_branchDest[0] .is_wysiwyg = "true";
defparam \temp_branchDest[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N15
dffeas \temp_branchDest[4] (
	.clk(CLK),
	.d(\temp_branchDest~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(ex_mem_flush3),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branchDest_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_branchDest[4] .is_wysiwyg = "true";
defparam \temp_branchDest[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N9
dffeas \temp_branchDest[3] (
	.clk(CLK),
	.d(\temp_branchDest~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(ex_mem_flush3),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branchDest_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_branchDest[3] .is_wysiwyg = "true";
defparam \temp_branchDest[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N7
dffeas \temp_branchDest[2] (
	.clk(CLK),
	.d(\temp_branchDest~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(ex_mem_flush3),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branchDest_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_branchDest[2] .is_wysiwyg = "true";
defparam \temp_branchDest[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N29
dffeas \temp_branchDest[1] (
	.clk(CLK),
	.d(\temp_branchDest~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(ex_mem_flush3),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branchDest_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_branchDest[1] .is_wysiwyg = "true";
defparam \temp_branchDest[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y42_N29
dffeas temp_zeroFlag(
	.clk(CLK),
	.d(Equal0),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(ex_mem_flush3),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_zeroFlag1),
	.prn(vcc));
// synopsys translate_off
defparam temp_zeroFlag.is_wysiwyg = "true";
defparam temp_zeroFlag.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N5
dffeas \temp_aluResult[1] (
	.clk(CLK),
	.d(\temp_aluResult~35_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[1] .is_wysiwyg = "true";
defparam \temp_aluResult[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N23
dffeas temp_dmemWEN(
	.clk(CLK),
	.d(\temp_dmemWEN~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dmemWEN1),
	.prn(vcc));
// synopsys translate_off
defparam temp_dmemWEN.is_wysiwyg = "true";
defparam temp_dmemWEN.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N13
dffeas temp_dmemREN(
	.clk(CLK),
	.d(\temp_dmemREN~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dmemREN1),
	.prn(vcc));
// synopsys translate_off
defparam temp_dmemREN.is_wysiwyg = "true";
defparam temp_dmemREN.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N15
dffeas \temp_aluResult[0] (
	.clk(CLK),
	.d(\temp_aluResult~36_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[0] .is_wysiwyg = "true";
defparam \temp_aluResult[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y42_N13
dffeas \temp_aluResult[2] (
	.clk(CLK),
	.d(\temp_aluResult~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[2] .is_wysiwyg = "true";
defparam \temp_aluResult[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N23
dffeas \temp_aluResult[3] (
	.clk(CLK),
	.d(\temp_aluResult~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[3] .is_wysiwyg = "true";
defparam \temp_aluResult[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N17
dffeas \temp_aluResult[5] (
	.clk(CLK),
	.d(\temp_aluResult~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[5] .is_wysiwyg = "true";
defparam \temp_aluResult[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N27
dffeas \temp_aluResult[4] (
	.clk(CLK),
	.d(\temp_aluResult~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[4] .is_wysiwyg = "true";
defparam \temp_aluResult[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N3
dffeas \temp_aluResult[7] (
	.clk(CLK),
	.d(\temp_aluResult~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[7] .is_wysiwyg = "true";
defparam \temp_aluResult[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N1
dffeas \temp_aluResult[6] (
	.clk(CLK),
	.d(\temp_aluResult~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[6] .is_wysiwyg = "true";
defparam \temp_aluResult[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N5
dffeas \temp_aluResult[9] (
	.clk(CLK),
	.d(\temp_aluResult~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[9] .is_wysiwyg = "true";
defparam \temp_aluResult[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N17
dffeas \temp_aluResult[8] (
	.clk(CLK),
	.d(\temp_aluResult~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[8] .is_wysiwyg = "true";
defparam \temp_aluResult[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y43_N13
dffeas \temp_aluResult[11] (
	.clk(CLK),
	.d(\temp_aluResult~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[11] .is_wysiwyg = "true";
defparam \temp_aluResult[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y43_N15
dffeas \temp_aluResult[10] (
	.clk(CLK),
	.d(\temp_aluResult~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[10] .is_wysiwyg = "true";
defparam \temp_aluResult[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N3
dffeas \temp_aluResult[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\temp_aluResult~15_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[13] .is_wysiwyg = "true";
defparam \temp_aluResult[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y43_N9
dffeas \temp_aluResult[12] (
	.clk(CLK),
	.d(\temp_aluResult~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[12] .is_wysiwyg = "true";
defparam \temp_aluResult[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N21
dffeas \temp_aluResult[15] (
	.clk(CLK),
	.d(\temp_aluResult~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[15] .is_wysiwyg = "true";
defparam \temp_aluResult[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y43_N1
dffeas \temp_aluResult[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\temp_aluResult~18_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[14] .is_wysiwyg = "true";
defparam \temp_aluResult[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y43_N23
dffeas \temp_aluResult[17] (
	.clk(CLK),
	.d(\temp_aluResult~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[17] .is_wysiwyg = "true";
defparam \temp_aluResult[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y43_N29
dffeas \temp_aluResult[16] (
	.clk(CLK),
	.d(\temp_aluResult~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[16] .is_wysiwyg = "true";
defparam \temp_aluResult[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y43_N7
dffeas \temp_aluResult[19] (
	.clk(CLK),
	.d(\temp_aluResult~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[19] .is_wysiwyg = "true";
defparam \temp_aluResult[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y43_N25
dffeas \temp_aluResult[18] (
	.clk(CLK),
	.d(\temp_aluResult~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[18] .is_wysiwyg = "true";
defparam \temp_aluResult[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y43_N27
dffeas \temp_aluResult[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\temp_aluResult~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[20] .is_wysiwyg = "true";
defparam \temp_aluResult[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N21
dffeas \temp_aluResult[21] (
	.clk(CLK),
	.d(\temp_aluResult~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[21] .is_wysiwyg = "true";
defparam \temp_aluResult[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N25
dffeas \temp_aluResult[23] (
	.clk(CLK),
	.d(\temp_aluResult~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[23] .is_wysiwyg = "true";
defparam \temp_aluResult[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N19
dffeas \temp_aluResult[22] (
	.clk(CLK),
	.d(\temp_aluResult~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[22] .is_wysiwyg = "true";
defparam \temp_aluResult[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N17
dffeas \temp_aluResult[25] (
	.clk(CLK),
	.d(\temp_aluResult~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[25] .is_wysiwyg = "true";
defparam \temp_aluResult[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N23
dffeas \temp_aluResult[24] (
	.clk(CLK),
	.d(\temp_aluResult~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[24] .is_wysiwyg = "true";
defparam \temp_aluResult[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N13
dffeas \temp_aluResult[26] (
	.clk(CLK),
	.d(\temp_aluResult~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[26] .is_wysiwyg = "true";
defparam \temp_aluResult[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N9
dffeas \temp_aluResult[27] (
	.clk(CLK),
	.d(\temp_aluResult~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[27] .is_wysiwyg = "true";
defparam \temp_aluResult[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N19
dffeas \temp_aluResult[29] (
	.clk(CLK),
	.d(\temp_aluResult~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[29] .is_wysiwyg = "true";
defparam \temp_aluResult[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N7
dffeas \temp_aluResult[28] (
	.clk(CLK),
	.d(\temp_aluResult~32_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[28] .is_wysiwyg = "true";
defparam \temp_aluResult[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N7
dffeas \temp_aluResult[31] (
	.clk(CLK),
	.d(\temp_aluResult~33_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[31] .is_wysiwyg = "true";
defparam \temp_aluResult[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N11
dffeas \temp_aluResult[30] (
	.clk(CLK),
	.d(\temp_aluResult~34_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[30] .is_wysiwyg = "true";
defparam \temp_aluResult[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y44_N13
dffeas temp_halt_out(
	.clk(CLK),
	.d(\temp_halt_out~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_halt_out1),
	.prn(vcc));
// synopsys translate_off
defparam temp_halt_out.is_wysiwyg = "true";
defparam temp_halt_out.power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N1
dffeas \temp_rdat2[0] (
	.clk(CLK),
	.d(\temp_rdat2~60_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[0] .is_wysiwyg = "true";
defparam \temp_rdat2[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N25
dffeas temp_regwrite(
	.clk(CLK),
	.d(\temp_regwrite~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_regwrite1),
	.prn(vcc));
// synopsys translate_off
defparam temp_regwrite.is_wysiwyg = "true";
defparam temp_regwrite.power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y44_N7
dffeas \temp_memtoreg[0] (
	.clk(CLK),
	.d(\temp_memtoreg~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_memtoreg_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_memtoreg[0] .is_wysiwyg = "true";
defparam \temp_memtoreg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N7
dffeas \temp_memtoreg[1] (
	.clk(CLK),
	.d(\temp_memtoreg~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_memtoreg_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_memtoreg[1] .is_wysiwyg = "true";
defparam \temp_memtoreg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N7
dffeas \temp_iMemLoad[0] (
	.clk(CLK),
	.d(\temp_iMemLoad~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[0] .is_wysiwyg = "true";
defparam \temp_iMemLoad[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N21
dffeas \temp_iMemLoad[15] (
	.clk(CLK),
	.d(\temp_iMemLoad~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[15] .is_wysiwyg = "true";
defparam \temp_iMemLoad[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y44_N23
dffeas \temp_iMemLoad[14] (
	.clk(CLK),
	.d(\temp_iMemLoad~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[14] .is_wysiwyg = "true";
defparam \temp_iMemLoad[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N5
dffeas \temp_iMemLoad[13] (
	.clk(CLK),
	.d(\temp_iMemLoad~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[13] .is_wysiwyg = "true";
defparam \temp_iMemLoad[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N5
dffeas \temp_iMemLoad[10] (
	.clk(CLK),
	.d(\temp_iMemLoad~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[10] .is_wysiwyg = "true";
defparam \temp_iMemLoad[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N19
dffeas \temp_iMemLoad[9] (
	.clk(CLK),
	.d(\temp_iMemLoad~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[9] .is_wysiwyg = "true";
defparam \temp_iMemLoad[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N5
dffeas \temp_iMemLoad[12] (
	.clk(CLK),
	.d(\temp_iMemLoad~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[12] .is_wysiwyg = "true";
defparam \temp_iMemLoad[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N31
dffeas \temp_iMemLoad[11] (
	.clk(CLK),
	.d(\temp_iMemLoad~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[11] .is_wysiwyg = "true";
defparam \temp_iMemLoad[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y42_N17
dffeas \temp_iMemLoad[1] (
	.clk(CLK),
	.d(\temp_iMemLoad~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[1] .is_wysiwyg = "true";
defparam \temp_iMemLoad[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y42_N27
dffeas \temp_iMemLoad[4] (
	.clk(CLK),
	.d(\temp_iMemLoad~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[4] .is_wysiwyg = "true";
defparam \temp_iMemLoad[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N31
dffeas \temp_iMemLoad[3] (
	.clk(CLK),
	.d(\temp_iMemLoad~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[3] .is_wysiwyg = "true";
defparam \temp_iMemLoad[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y44_N17
dffeas \temp_iMemLoad[2] (
	.clk(CLK),
	.d(\temp_iMemLoad~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[2] .is_wysiwyg = "true";
defparam \temp_iMemLoad[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N5
dffeas \temp_iMemLoad[8] (
	.clk(CLK),
	.d(\temp_iMemLoad~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[8] .is_wysiwyg = "true";
defparam \temp_iMemLoad[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N19
dffeas \temp_iMemLoad[7] (
	.clk(CLK),
	.d(\temp_iMemLoad~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[7] .is_wysiwyg = "true";
defparam \temp_iMemLoad[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N25
dffeas \temp_iMemLoad[6] (
	.clk(CLK),
	.d(\temp_iMemLoad~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[6] .is_wysiwyg = "true";
defparam \temp_iMemLoad[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N23
dffeas \temp_iMemLoad[5] (
	.clk(CLK),
	.d(\temp_iMemLoad~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[5] .is_wysiwyg = "true";
defparam \temp_iMemLoad[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N7
dffeas \temp_iMemLoad[31] (
	.clk(CLK),
	.d(\temp_iMemLoad~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[31] .is_wysiwyg = "true";
defparam \temp_iMemLoad[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N29
dffeas \temp_iMemLoad[30] (
	.clk(CLK),
	.d(\temp_iMemLoad~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[30] .is_wysiwyg = "true";
defparam \temp_iMemLoad[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N25
dffeas \temp_iMemLoad[29] (
	.clk(CLK),
	.d(\temp_iMemLoad~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[29] .is_wysiwyg = "true";
defparam \temp_iMemLoad[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y42_N1
dffeas \temp_iMemLoad[27] (
	.clk(CLK),
	.d(\temp_iMemLoad~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[27] .is_wysiwyg = "true";
defparam \temp_iMemLoad[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y42_N19
dffeas \temp_iMemLoad[26] (
	.clk(CLK),
	.d(\temp_iMemLoad~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[26] .is_wysiwyg = "true";
defparam \temp_iMemLoad[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y42_N29
dffeas \temp_iMemLoad[28] (
	.clk(CLK),
	.d(\temp_iMemLoad~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[28] .is_wysiwyg = "true";
defparam \temp_iMemLoad[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N3
dffeas temp_branchSelect(
	.clk(CLK),
	.d(\temp_branchSelect~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branchSelect1),
	.prn(vcc));
// synopsys translate_off
defparam temp_branchSelect.is_wysiwyg = "true";
defparam temp_branchSelect.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y42_N31
dffeas \temp_rdat1[1] (
	.clk(CLK),
	.d(\temp_rdat1~63_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[1] .is_wysiwyg = "true";
defparam \temp_rdat1[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N15
dffeas \temp_npc[1] (
	.clk(CLK),
	.d(\temp_npc~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[1] .is_wysiwyg = "true";
defparam \temp_npc[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N1
dffeas \temp_pcselect[1] (
	.clk(CLK),
	.d(\temp_pcselect~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_pcselect_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_pcselect[1] .is_wysiwyg = "true";
defparam \temp_pcselect[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y42_N17
dffeas \temp_pcselect[0] (
	.clk(CLK),
	.d(\temp_pcselect~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_pcselect_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_pcselect[0] .is_wysiwyg = "true";
defparam \temp_pcselect[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y42_N9
dffeas \temp_rdat1[0] (
	.clk(CLK),
	.d(\temp_rdat1~64_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[0] .is_wysiwyg = "true";
defparam \temp_rdat1[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N29
dffeas \temp_npc[0] (
	.clk(CLK),
	.d(\temp_npc~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[0] .is_wysiwyg = "true";
defparam \temp_npc[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N19
dffeas \temp_npc[2] (
	.clk(CLK),
	.d(\temp_npc~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[2] .is_wysiwyg = "true";
defparam \temp_npc[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N25
dffeas \temp_rdat1[2] (
	.clk(CLK),
	.d(\temp_rdat1~65_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[2] .is_wysiwyg = "true";
defparam \temp_rdat1[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N11
dffeas \temp_npc[3] (
	.clk(CLK),
	.d(\temp_npc~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[3] .is_wysiwyg = "true";
defparam \temp_npc[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N23
dffeas \temp_rdat1[3] (
	.clk(CLK),
	.d(\temp_rdat1~62_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[3] .is_wysiwyg = "true";
defparam \temp_rdat1[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N15
dffeas \temp_npc[5] (
	.clk(CLK),
	.d(\temp_npc~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[5] .is_wysiwyg = "true";
defparam \temp_npc[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y44_N1
dffeas \temp_npc[4] (
	.clk(CLK),
	.d(\temp_npc~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[4] .is_wysiwyg = "true";
defparam \temp_npc[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N29
dffeas \temp_rdat1[5] (
	.clk(CLK),
	.d(\temp_rdat1~66_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[5] .is_wysiwyg = "true";
defparam \temp_rdat1[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y44_N11
dffeas \temp_rdat1[4] (
	.clk(CLK),
	.d(\temp_rdat1~67_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[4] .is_wysiwyg = "true";
defparam \temp_rdat1[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N3
dffeas \temp_npc[7] (
	.clk(CLK),
	.d(\temp_npc~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[7] .is_wysiwyg = "true";
defparam \temp_npc[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N21
dffeas \temp_npc[6] (
	.clk(CLK),
	.d(\temp_npc~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[6] .is_wysiwyg = "true";
defparam \temp_npc[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N25
dffeas \temp_rdat1[7] (
	.clk(CLK),
	.d(\temp_rdat1~68_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[7] .is_wysiwyg = "true";
defparam \temp_rdat1[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y45_N1
dffeas \temp_rdat1[6] (
	.clk(CLK),
	.d(\temp_rdat1[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[6] .is_wysiwyg = "true";
defparam \temp_rdat1[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N9
dffeas \temp_npc[9] (
	.clk(CLK),
	.d(\temp_npc~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[9] .is_wysiwyg = "true";
defparam \temp_npc[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N29
dffeas \temp_npc[8] (
	.clk(CLK),
	.d(\temp_npc~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[8] .is_wysiwyg = "true";
defparam \temp_npc[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N7
dffeas \temp_rdat1[9] (
	.clk(CLK),
	.d(\temp_rdat1~70_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[9] .is_wysiwyg = "true";
defparam \temp_rdat1[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y45_N7
dffeas \temp_rdat1[8] (
	.clk(CLK),
	.d(\temp_rdat1~71_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[8] .is_wysiwyg = "true";
defparam \temp_rdat1[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N19
dffeas \temp_npc[11] (
	.clk(CLK),
	.d(\temp_npc~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[11] .is_wysiwyg = "true";
defparam \temp_npc[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N19
dffeas \temp_npc[10] (
	.clk(CLK),
	.d(\temp_npc~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[10] .is_wysiwyg = "true";
defparam \temp_npc[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N1
dffeas \temp_rdat1[11] (
	.clk(CLK),
	.d(\temp_rdat1~72_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[11] .is_wysiwyg = "true";
defparam \temp_rdat1[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y45_N17
dffeas \temp_rdat1[10] (
	.clk(CLK),
	.d(\temp_rdat1~73_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[10] .is_wysiwyg = "true";
defparam \temp_rdat1[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N1
dffeas \temp_npc[13] (
	.clk(CLK),
	.d(\temp_npc~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[13] .is_wysiwyg = "true";
defparam \temp_npc[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N9
dffeas \temp_npc[12] (
	.clk(CLK),
	.d(\temp_npc~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[12] .is_wysiwyg = "true";
defparam \temp_npc[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N17
dffeas \temp_rdat1[13] (
	.clk(CLK),
	.d(\temp_rdat1~74_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[13] .is_wysiwyg = "true";
defparam \temp_rdat1[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y45_N27
dffeas \temp_rdat1[12] (
	.clk(CLK),
	.d(\temp_rdat1~75_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[12] .is_wysiwyg = "true";
defparam \temp_rdat1[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N25
dffeas \temp_npc[15] (
	.clk(CLK),
	.d(\temp_npc~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[15] .is_wysiwyg = "true";
defparam \temp_npc[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N23
dffeas \temp_npc[14] (
	.clk(CLK),
	.d(\temp_npc~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[14] .is_wysiwyg = "true";
defparam \temp_npc[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N13
dffeas \temp_rdat1[15] (
	.clk(CLK),
	.d(\temp_rdat1~76_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[15] .is_wysiwyg = "true";
defparam \temp_rdat1[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N3
dffeas \temp_rdat1[14] (
	.clk(CLK),
	.d(\temp_rdat1~77_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[14] .is_wysiwyg = "true";
defparam \temp_rdat1[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N21
dffeas \temp_npc[17] (
	.clk(CLK),
	.d(\temp_npc~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[17] .is_wysiwyg = "true";
defparam \temp_npc[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N3
dffeas \temp_npc[16] (
	.clk(CLK),
	.d(\temp_npc~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[16] .is_wysiwyg = "true";
defparam \temp_npc[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N9
dffeas \temp_rdat1[17] (
	.clk(CLK),
	.d(\temp_rdat1~78_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[17] .is_wysiwyg = "true";
defparam \temp_rdat1[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y44_N9
dffeas \temp_rdat1[16] (
	.clk(CLK),
	.d(\temp_rdat1~79_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[16] .is_wysiwyg = "true";
defparam \temp_rdat1[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N3
dffeas \temp_signZero[16] (
	.clk(CLK),
	.d(\temp_signZero~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_signZero_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_signZero[16] .is_wysiwyg = "true";
defparam \temp_signZero[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N29
dffeas \temp_npc[19] (
	.clk(CLK),
	.d(\temp_npc~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[19] .is_wysiwyg = "true";
defparam \temp_npc[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N5
dffeas \temp_npc[18] (
	.clk(CLK),
	.d(\temp_npc~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[18] .is_wysiwyg = "true";
defparam \temp_npc[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N1
dffeas \temp_rdat1[19] (
	.clk(CLK),
	.d(\temp_rdat1~80_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[19] .is_wysiwyg = "true";
defparam \temp_rdat1[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y45_N1
dffeas \temp_iMemLoad[17] (
	.clk(CLK),
	.d(\temp_iMemLoad~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[17] .is_wysiwyg = "true";
defparam \temp_iMemLoad[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N15
dffeas \temp_rdat1[18] (
	.clk(CLK),
	.d(\temp_rdat1~81_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[18] .is_wysiwyg = "true";
defparam \temp_rdat1[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N15
dffeas \temp_iMemLoad[16] (
	.clk(CLK),
	.d(\temp_iMemLoad~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[16] .is_wysiwyg = "true";
defparam \temp_iMemLoad[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N7
dffeas \temp_npc[20] (
	.clk(CLK),
	.d(\temp_npc~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[20] .is_wysiwyg = "true";
defparam \temp_npc[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y45_N27
dffeas \temp_rdat1[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\temp_rdat1~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[20] .is_wysiwyg = "true";
defparam \temp_rdat1[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y44_N1
dffeas \temp_iMemLoad[18] (
	.clk(CLK),
	.d(\temp_iMemLoad~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[18] .is_wysiwyg = "true";
defparam \temp_iMemLoad[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N13
dffeas \temp_npc[21] (
	.clk(CLK),
	.d(\temp_npc~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[21] .is_wysiwyg = "true";
defparam \temp_npc[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N9
dffeas \temp_rdat1[21] (
	.clk(CLK),
	.d(\temp_rdat1~83_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[21] .is_wysiwyg = "true";
defparam \temp_rdat1[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N5
dffeas \temp_iMemLoad[19] (
	.clk(CLK),
	.d(\temp_iMemLoad~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[19] .is_wysiwyg = "true";
defparam \temp_iMemLoad[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N3
dffeas \temp_npc[23] (
	.clk(CLK),
	.d(\temp_npc~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[23] .is_wysiwyg = "true";
defparam \temp_npc[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y44_N31
dffeas \temp_npc[22] (
	.clk(CLK),
	.d(\temp_npc~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[22] .is_wysiwyg = "true";
defparam \temp_npc[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y44_N19
dffeas \temp_rdat1[23] (
	.clk(CLK),
	.d(\temp_rdat1~84_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[23] .is_wysiwyg = "true";
defparam \temp_rdat1[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y44_N3
dffeas \temp_iMemLoad[21] (
	.clk(CLK),
	.d(\temp_iMemLoad~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[21] .is_wysiwyg = "true";
defparam \temp_iMemLoad[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y44_N3
dffeas \temp_rdat1[22] (
	.clk(CLK),
	.d(\temp_rdat1~85_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[22] .is_wysiwyg = "true";
defparam \temp_rdat1[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y44_N11
dffeas \temp_iMemLoad[20] (
	.clk(CLK),
	.d(\temp_iMemLoad~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[20] .is_wysiwyg = "true";
defparam \temp_iMemLoad[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N13
dffeas \temp_npc[25] (
	.clk(CLK),
	.d(\temp_npc~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[25] .is_wysiwyg = "true";
defparam \temp_npc[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y44_N11
dffeas \temp_npc[24] (
	.clk(CLK),
	.d(\temp_npc~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[24] .is_wysiwyg = "true";
defparam \temp_npc[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N1
dffeas \temp_rdat1[25] (
	.clk(CLK),
	.d(\temp_rdat1~86_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[25] .is_wysiwyg = "true";
defparam \temp_rdat1[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N15
dffeas \temp_iMemLoad[23] (
	.clk(CLK),
	.d(\temp_iMemLoad~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[23] .is_wysiwyg = "true";
defparam \temp_iMemLoad[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y44_N17
dffeas \temp_rdat1[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\temp_rdat1~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[24] .is_wysiwyg = "true";
defparam \temp_rdat1[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y44_N31
dffeas \temp_iMemLoad[22] (
	.clk(CLK),
	.d(\temp_iMemLoad~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_iMemLoad_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_iMemLoad[22] .is_wysiwyg = "true";
defparam \temp_iMemLoad[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N3
dffeas \temp_npc[26] (
	.clk(CLK),
	.d(\temp_npc~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[26] .is_wysiwyg = "true";
defparam \temp_npc[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N9
dffeas \temp_rdat1[26] (
	.clk(CLK),
	.d(\temp_rdat1~88_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[26] .is_wysiwyg = "true";
defparam \temp_rdat1[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N5
dffeas \temp_npc[27] (
	.clk(CLK),
	.d(\temp_npc~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[27] .is_wysiwyg = "true";
defparam \temp_npc[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y44_N19
dffeas \temp_rdat1[27] (
	.clk(CLK),
	.d(\temp_rdat1~89_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[27] .is_wysiwyg = "true";
defparam \temp_rdat1[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N19
dffeas \temp_npc[29] (
	.clk(CLK),
	.d(\temp_npc~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[29] .is_wysiwyg = "true";
defparam \temp_npc[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N11
dffeas \temp_npc[28] (
	.clk(CLK),
	.d(\temp_npc~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[28] .is_wysiwyg = "true";
defparam \temp_npc[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y44_N23
dffeas \temp_rdat1[29] (
	.clk(CLK),
	.d(\temp_rdat1~90_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[29] .is_wysiwyg = "true";
defparam \temp_rdat1[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y44_N13
dffeas \temp_rdat1[28] (
	.clk(CLK),
	.d(\temp_rdat1~91_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[28] .is_wysiwyg = "true";
defparam \temp_rdat1[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N19
dffeas \temp_rdat1[31] (
	.clk(CLK),
	.d(\temp_rdat1~92_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[31] .is_wysiwyg = "true";
defparam \temp_rdat1[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y44_N31
dffeas \temp_npc[31] (
	.clk(CLK),
	.d(\temp_npc~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[31] .is_wysiwyg = "true";
defparam \temp_npc[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N13
dffeas \temp_npc[30] (
	.clk(CLK),
	.d(\temp_npc~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[30] .is_wysiwyg = "true";
defparam \temp_npc[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y42_N13
dffeas \temp_rdat1[30] (
	.clk(CLK),
	.d(\temp_rdat1~93_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat1_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat1[30] .is_wysiwyg = "true";
defparam \temp_rdat1[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N7
dffeas \temp_rdat2[1] (
	.clk(CLK),
	.d(\temp_rdat2~61_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[1] .is_wysiwyg = "true";
defparam \temp_rdat2[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N29
dffeas \temp_rdat2[2] (
	.clk(CLK),
	.d(\temp_rdat2~62_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[2] .is_wysiwyg = "true";
defparam \temp_rdat2[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N5
dffeas \temp_rdat2[3] (
	.clk(CLK),
	.d(\temp_rdat2~63_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[3] .is_wysiwyg = "true";
defparam \temp_rdat2[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N17
dffeas \temp_rdat2[4] (
	.clk(CLK),
	.d(\temp_rdat2~64_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[4] .is_wysiwyg = "true";
defparam \temp_rdat2[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N15
dffeas \temp_rdat2[5] (
	.clk(CLK),
	.d(\temp_rdat2~65_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[5] .is_wysiwyg = "true";
defparam \temp_rdat2[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y42_N31
dffeas \temp_rdat2[6] (
	.clk(CLK),
	.d(\temp_rdat2~66_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[6] .is_wysiwyg = "true";
defparam \temp_rdat2[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N15
dffeas \temp_rdat2[7] (
	.clk(CLK),
	.d(\temp_rdat2~67_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[7] .is_wysiwyg = "true";
defparam \temp_rdat2[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N11
dffeas \temp_rdat2[8] (
	.clk(CLK),
	.d(\temp_rdat2~68_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[8] .is_wysiwyg = "true";
defparam \temp_rdat2[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N21
dffeas \temp_rdat2[9] (
	.clk(CLK),
	.d(\temp_rdat2~69_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[9] .is_wysiwyg = "true";
defparam \temp_rdat2[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N9
dffeas \temp_rdat2[10] (
	.clk(CLK),
	.d(\temp_rdat2~70_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[10] .is_wysiwyg = "true";
defparam \temp_rdat2[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y44_N25
dffeas \temp_rdat2[11] (
	.clk(CLK),
	.d(\temp_rdat2~71_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[11] .is_wysiwyg = "true";
defparam \temp_rdat2[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N3
dffeas \temp_rdat2[12] (
	.clk(CLK),
	.d(\temp_rdat2~72_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[12] .is_wysiwyg = "true";
defparam \temp_rdat2[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N27
dffeas \temp_rdat2[13] (
	.clk(CLK),
	.d(\temp_rdat2~73_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[13] .is_wysiwyg = "true";
defparam \temp_rdat2[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N21
dffeas \temp_rdat2[14] (
	.clk(CLK),
	.d(\temp_rdat2~74_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[14] .is_wysiwyg = "true";
defparam \temp_rdat2[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y37_N27
dffeas \temp_rdat2[15] (
	.clk(CLK),
	.d(\temp_rdat2~75_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[15] .is_wysiwyg = "true";
defparam \temp_rdat2[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N31
dffeas \temp_rdat2[16] (
	.clk(CLK),
	.d(\temp_rdat2~76_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[16] .is_wysiwyg = "true";
defparam \temp_rdat2[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N19
dffeas \temp_rdat2[17] (
	.clk(CLK),
	.d(\temp_rdat2~77_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[17] .is_wysiwyg = "true";
defparam \temp_rdat2[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y37_N25
dffeas \temp_rdat2[18] (
	.clk(CLK),
	.d(\temp_rdat2~78_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[18] .is_wysiwyg = "true";
defparam \temp_rdat2[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y37_N31
dffeas \temp_rdat2[19] (
	.clk(CLK),
	.d(\temp_rdat2~79_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[19] .is_wysiwyg = "true";
defparam \temp_rdat2[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N9
dffeas \temp_rdat2[20] (
	.clk(CLK),
	.d(\temp_rdat2~80_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[20] .is_wysiwyg = "true";
defparam \temp_rdat2[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N27
dffeas \temp_rdat2[21] (
	.clk(CLK),
	.d(\temp_rdat2~81_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[21] .is_wysiwyg = "true";
defparam \temp_rdat2[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y42_N27
dffeas \temp_rdat2[22] (
	.clk(CLK),
	.d(\temp_rdat2~82_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[22] .is_wysiwyg = "true";
defparam \temp_rdat2[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N25
dffeas \temp_rdat2[23] (
	.clk(CLK),
	.d(\temp_rdat2~83_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[23] .is_wysiwyg = "true";
defparam \temp_rdat2[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N25
dffeas \temp_rdat2[24] (
	.clk(CLK),
	.d(\temp_rdat2~84_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[24] .is_wysiwyg = "true";
defparam \temp_rdat2[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N11
dffeas \temp_rdat2[25] (
	.clk(CLK),
	.d(\temp_rdat2~85_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[25] .is_wysiwyg = "true";
defparam \temp_rdat2[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N23
dffeas \temp_rdat2[26] (
	.clk(CLK),
	.d(\temp_rdat2~86_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[26] .is_wysiwyg = "true";
defparam \temp_rdat2[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y37_N29
dffeas \temp_rdat2[27] (
	.clk(CLK),
	.d(\temp_rdat2~87_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[27] .is_wysiwyg = "true";
defparam \temp_rdat2[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N17
dffeas \temp_rdat2[28] (
	.clk(CLK),
	.d(\temp_rdat2~88_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[28] .is_wysiwyg = "true";
defparam \temp_rdat2[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N15
dffeas \temp_rdat2[29] (
	.clk(CLK),
	.d(\temp_rdat2~89_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[29] .is_wysiwyg = "true";
defparam \temp_rdat2[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y37_N19
dffeas \temp_rdat2[30] (
	.clk(CLK),
	.d(\temp_rdat2~90_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[30] .is_wysiwyg = "true";
defparam \temp_rdat2[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N7
dffeas \temp_rdat2[31] (
	.clk(CLK),
	.d(\temp_rdat2~91_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat2_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat2[31] .is_wysiwyg = "true";
defparam \temp_rdat2[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N4
cycloneive_lcell_comb \temp_branchDest~0 (
// Equation(s):
// \temp_branchDest~0_combout  = (temp_regdst_output_0 & (((temp_imemload_output_11)))) # (!temp_regdst_output_0 & ((temp_regdst_output_1) # ((temp_imemload_output_16))))

	.dataa(temp_regdst_output_0),
	.datab(temp_regdst_output_1),
	.datac(temp_imemload_output_16),
	.datad(temp_imemload_output_11),
	.cin(gnd),
	.combout(\temp_branchDest~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_branchDest~0 .lut_mask = 16'hFE54;
defparam \temp_branchDest~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N14
cycloneive_lcell_comb \temp_branchDest~1 (
// Equation(s):
// \temp_branchDest~1_combout  = (temp_regdst_output_0 & (((temp_imemload_output_15)))) # (!temp_regdst_output_0 & ((temp_regdst_output_1) # ((temp_imemload_output_20))))

	.dataa(temp_regdst_output_0),
	.datab(temp_regdst_output_1),
	.datac(temp_imemload_output_15),
	.datad(temp_imemload_output_20),
	.cin(gnd),
	.combout(\temp_branchDest~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_branchDest~1 .lut_mask = 16'hF5E4;
defparam \temp_branchDest~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N8
cycloneive_lcell_comb \temp_branchDest~2 (
// Equation(s):
// \temp_branchDest~2_combout  = (temp_regdst_output_0 & (((temp_imemload_output_14)))) # (!temp_regdst_output_0 & ((temp_imemload_output_19) # ((temp_regdst_output_1))))

	.dataa(temp_regdst_output_0),
	.datab(temp_imemload_output_19),
	.datac(temp_imemload_output_14),
	.datad(temp_regdst_output_1),
	.cin(gnd),
	.combout(\temp_branchDest~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_branchDest~2 .lut_mask = 16'hF5E4;
defparam \temp_branchDest~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N6
cycloneive_lcell_comb \temp_branchDest~3 (
// Equation(s):
// \temp_branchDest~3_combout  = (temp_regdst_output_0 & (((temp_imemload_output_13)))) # (!temp_regdst_output_0 & ((temp_regdst_output_1) # ((temp_imemload_output_18))))

	.dataa(temp_regdst_output_0),
	.datab(temp_regdst_output_1),
	.datac(temp_imemload_output_13),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\temp_branchDest~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_branchDest~3 .lut_mask = 16'hF5E4;
defparam \temp_branchDest~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N28
cycloneive_lcell_comb \temp_branchDest~4 (
// Equation(s):
// \temp_branchDest~4_combout  = (temp_regdst_output_0 & (((temp_imemload_output_12)))) # (!temp_regdst_output_0 & ((temp_imemload_output_17) # ((temp_regdst_output_1))))

	.dataa(temp_regdst_output_0),
	.datab(temp_imemload_output_17),
	.datac(temp_imemload_output_12),
	.datad(temp_regdst_output_1),
	.cin(gnd),
	.combout(\temp_branchDest~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_branchDest~4 .lut_mask = 16'hF5E4;
defparam \temp_branchDest~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N4
cycloneive_lcell_comb \temp_aluResult~35 (
// Equation(s):
// \temp_aluResult~35_combout  = (Mux302 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(Mux30),
	.cin(gnd),
	.combout(\temp_aluResult~35_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~35 .lut_mask = 16'h5700;
defparam \temp_aluResult~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N26
cycloneive_lcell_comb \temp_dmemWEN~0 (
// Equation(s):
// \temp_dmemWEN~0_combout  = (temp_request_dmemWEN_output1 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(temp_request_dmemWEN_output),
	.cin(gnd),
	.combout(\temp_dmemWEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dmemWEN~0 .lut_mask = 16'h1F00;
defparam \temp_dmemWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N22
cycloneive_lcell_comb \temp_dmemWEN~feeder (
// Equation(s):
// \temp_dmemWEN~feeder_combout  = \temp_dmemWEN~0_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\temp_dmemWEN~0_combout ),
	.cin(gnd),
	.combout(\temp_dmemWEN~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dmemWEN~feeder .lut_mask = 16'hFF00;
defparam \temp_dmemWEN~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N30
cycloneive_lcell_comb \temp_dmemREN~0 (
// Equation(s):
// \temp_dmemREN~0_combout  = (temp_request_dmemREN_output1 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(temp_request_dmemREN_output),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_dmemREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dmemREN~0 .lut_mask = 16'h04CC;
defparam \temp_dmemREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N12
cycloneive_lcell_comb \temp_dmemREN~feeder (
// Equation(s):
// \temp_dmemREN~feeder_combout  = \temp_dmemREN~0_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\temp_dmemREN~0_combout ),
	.cin(gnd),
	.combout(\temp_dmemREN~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dmemREN~feeder .lut_mask = 16'hFF00;
defparam \temp_dmemREN~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N14
cycloneive_lcell_comb \temp_aluResult~36 (
// Equation(s):
// \temp_aluResult~36_combout  = (Mux312 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(Mux31),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_aluResult~36_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~36 .lut_mask = 16'h10F0;
defparam \temp_aluResult~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N12
cycloneive_lcell_comb \temp_aluResult~4 (
// Equation(s):
// \temp_aluResult~4_combout  = (!ex_mem_flush3 & (!temp_ALUop_output_3 & Mux292))

	.dataa(ex_mem_flush3),
	.datab(gnd),
	.datac(temp_ALUop_output_3),
	.datad(Mux29),
	.cin(gnd),
	.combout(\temp_aluResult~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~4 .lut_mask = 16'h0500;
defparam \temp_aluResult~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N22
cycloneive_lcell_comb \temp_aluResult~5 (
// Equation(s):
// \temp_aluResult~5_combout  = (!ex_mem_flush3 & (!temp_ALUop_output_3 & Mux282))

	.dataa(ex_mem_flush3),
	.datab(gnd),
	.datac(temp_ALUop_output_3),
	.datad(Mux28),
	.cin(gnd),
	.combout(\temp_aluResult~5_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~5 .lut_mask = 16'h0500;
defparam \temp_aluResult~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N16
cycloneive_lcell_comb \temp_aluResult~6 (
// Equation(s):
// \temp_aluResult~6_combout  = (!temp_ALUop_output_3 & (!ex_mem_flush3 & Mux261))

	.dataa(gnd),
	.datab(temp_ALUop_output_3),
	.datac(ex_mem_flush3),
	.datad(Mux26),
	.cin(gnd),
	.combout(\temp_aluResult~6_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~6 .lut_mask = 16'h0300;
defparam \temp_aluResult~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N26
cycloneive_lcell_comb \temp_aluResult~7 (
// Equation(s):
// \temp_aluResult~7_combout  = (!ex_mem_flush3 & (Mux272 & !temp_ALUop_output_3))

	.dataa(ex_mem_flush3),
	.datab(Mux27),
	.datac(gnd),
	.datad(temp_ALUop_output_3),
	.cin(gnd),
	.combout(\temp_aluResult~7_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~7 .lut_mask = 16'h0044;
defparam \temp_aluResult~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N2
cycloneive_lcell_comb \temp_aluResult~8 (
// Equation(s):
// \temp_aluResult~8_combout  = (!temp_ALUop_output_3 & (!ex_mem_flush3 & Mux241))

	.dataa(temp_ALUop_output_3),
	.datab(gnd),
	.datac(ex_mem_flush3),
	.datad(Mux24),
	.cin(gnd),
	.combout(\temp_aluResult~8_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~8 .lut_mask = 16'h0500;
defparam \temp_aluResult~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N0
cycloneive_lcell_comb \temp_aluResult~9 (
// Equation(s):
// \temp_aluResult~9_combout  = (!temp_ALUop_output_3 & (!ex_mem_flush3 & Mux251))

	.dataa(temp_ALUop_output_3),
	.datab(gnd),
	.datac(ex_mem_flush3),
	.datad(Mux25),
	.cin(gnd),
	.combout(\temp_aluResult~9_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~9 .lut_mask = 16'h0500;
defparam \temp_aluResult~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N8
cycloneive_lcell_comb \temp_aluResult~10 (
// Equation(s):
// \temp_aluResult~10_combout  = (temp_ALUop_output_3) # ((ex_mem_flush & ((ex_mem_flush2) # (ex_mem_flush1))))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(temp_ALUop_output_3),
	.cin(gnd),
	.combout(\temp_aluResult~10_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~10 .lut_mask = 16'hFFE0;
defparam \temp_aluResult~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N4
cycloneive_lcell_comb \temp_aluResult~11 (
// Equation(s):
// \temp_aluResult~11_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & ((Mux221))) # (!Mux191 & (Mux222))))

	.dataa(Mux221),
	.datab(Mux22),
	.datac(\temp_aluResult~10_combout ),
	.datad(Mux19),
	.cin(gnd),
	.combout(\temp_aluResult~11_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~11 .lut_mask = 16'h0C0A;
defparam \temp_aluResult~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N16
cycloneive_lcell_comb \temp_aluResult~12 (
// Equation(s):
// \temp_aluResult~12_combout  = (!\temp_aluResult~10_combout  & ((Mux231) # ((!Mux191 & Mux232))))

	.dataa(Mux23),
	.datab(Mux19),
	.datac(\temp_aluResult~10_combout ),
	.datad(Mux231),
	.cin(gnd),
	.combout(\temp_aluResult~12_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~12 .lut_mask = 16'h0B0A;
defparam \temp_aluResult~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N12
cycloneive_lcell_comb \temp_aluResult~13 (
// Equation(s):
// \temp_aluResult~13_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux201)) # (!Mux191 & ((Mux202)))))

	.dataa(Mux19),
	.datab(Mux20),
	.datac(Mux201),
	.datad(\temp_aluResult~10_combout ),
	.cin(gnd),
	.combout(\temp_aluResult~13_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~13 .lut_mask = 16'h00D8;
defparam \temp_aluResult~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N14
cycloneive_lcell_comb \temp_aluResult~14 (
// Equation(s):
// \temp_aluResult~14_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux211)) # (!Mux191 & ((Mux212)))))

	.dataa(Mux19),
	.datab(Mux21),
	.datac(Mux211),
	.datad(\temp_aluResult~10_combout ),
	.cin(gnd),
	.combout(\temp_aluResult~14_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~14 .lut_mask = 16'h00D8;
defparam \temp_aluResult~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N0
cycloneive_lcell_comb \temp_aluResult~15 (
// Equation(s):
// \temp_aluResult~15_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux181)) # (!Mux191 & ((Mux182)))))

	.dataa(Mux19),
	.datab(Mux18),
	.datac(\temp_aluResult~10_combout ),
	.datad(Mux181),
	.cin(gnd),
	.combout(\temp_aluResult~15_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~15 .lut_mask = 16'h0D08;
defparam \temp_aluResult~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N8
cycloneive_lcell_comb \temp_aluResult~16 (
// Equation(s):
// \temp_aluResult~16_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & ((Mux192))) # (!Mux191 & (Mux193))))

	.dataa(\temp_aluResult~10_combout ),
	.datab(Mux19),
	.datac(Mux192),
	.datad(Mux191),
	.cin(gnd),
	.combout(\temp_aluResult~16_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~16 .lut_mask = 16'h5410;
defparam \temp_aluResult~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N20
cycloneive_lcell_comb \temp_aluResult~17 (
// Equation(s):
// \temp_aluResult~17_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux162)) # (!Mux191 & ((Mux163)))))

	.dataa(Mux16),
	.datab(Mux19),
	.datac(\temp_aluResult~10_combout ),
	.datad(Mux161),
	.cin(gnd),
	.combout(\temp_aluResult~17_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~17 .lut_mask = 16'h0B08;
defparam \temp_aluResult~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N20
cycloneive_lcell_comb \temp_aluResult~18 (
// Equation(s):
// \temp_aluResult~18_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux172)) # (!Mux191 & ((Mux173)))))

	.dataa(Mux17),
	.datab(Mux19),
	.datac(Mux171),
	.datad(\temp_aluResult~10_combout ),
	.cin(gnd),
	.combout(\temp_aluResult~18_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~18 .lut_mask = 16'h00B8;
defparam \temp_aluResult~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N22
cycloneive_lcell_comb \temp_aluResult~19 (
// Equation(s):
// \temp_aluResult~19_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux141)) # (!Mux191 & ((Mux142)))))

	.dataa(\temp_aluResult~10_combout ),
	.datab(Mux14),
	.datac(Mux141),
	.datad(Mux19),
	.cin(gnd),
	.combout(\temp_aluResult~19_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~19 .lut_mask = 16'h4450;
defparam \temp_aluResult~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N28
cycloneive_lcell_comb \temp_aluResult~20 (
// Equation(s):
// \temp_aluResult~20_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux151)) # (!Mux191 & ((Mux152)))))

	.dataa(Mux19),
	.datab(Mux15),
	.datac(Mux151),
	.datad(\temp_aluResult~10_combout ),
	.cin(gnd),
	.combout(\temp_aluResult~20_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~20 .lut_mask = 16'h00D8;
defparam \temp_aluResult~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N6
cycloneive_lcell_comb \temp_aluResult~21 (
// Equation(s):
// \temp_aluResult~21_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & ((Mux121))) # (!Mux191 & (Mux122))))

	.dataa(\temp_aluResult~10_combout ),
	.datab(Mux121),
	.datac(Mux19),
	.datad(Mux12),
	.cin(gnd),
	.combout(\temp_aluResult~21_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~21 .lut_mask = 16'h5404;
defparam \temp_aluResult~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N24
cycloneive_lcell_comb \temp_aluResult~22 (
// Equation(s):
// \temp_aluResult~22_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux131)) # (!Mux191 & ((Mux132)))))

	.dataa(Mux19),
	.datab(Mux13),
	.datac(\temp_aluResult~10_combout ),
	.datad(Mux131),
	.cin(gnd),
	.combout(\temp_aluResult~22_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~22 .lut_mask = 16'h0D08;
defparam \temp_aluResult~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N0
cycloneive_lcell_comb \temp_aluResult~23 (
// Equation(s):
// \temp_aluResult~23_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux111)) # (!Mux191 & ((Mux112)))))

	.dataa(\temp_aluResult~10_combout ),
	.datab(Mux19),
	.datac(Mux11),
	.datad(Mux111),
	.cin(gnd),
	.combout(\temp_aluResult~23_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~23 .lut_mask = 16'h5140;
defparam \temp_aluResult~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N20
cycloneive_lcell_comb \temp_aluResult~24 (
// Equation(s):
// \temp_aluResult~24_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux101)) # (!Mux191 & ((Mux102)))))

	.dataa(Mux10),
	.datab(Mux19),
	.datac(\temp_aluResult~10_combout ),
	.datad(Mux101),
	.cin(gnd),
	.combout(\temp_aluResult~24_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~24 .lut_mask = 16'h0B08;
defparam \temp_aluResult~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N24
cycloneive_lcell_comb \temp_aluResult~25 (
// Equation(s):
// \temp_aluResult~25_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux81)) # (!Mux191 & ((Mux82)))))

	.dataa(Mux8),
	.datab(\temp_aluResult~10_combout ),
	.datac(Mux19),
	.datad(Mux81),
	.cin(gnd),
	.combout(\temp_aluResult~25_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~25 .lut_mask = 16'h2320;
defparam \temp_aluResult~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N18
cycloneive_lcell_comb \temp_aluResult~26 (
// Equation(s):
// \temp_aluResult~26_combout  = (!\temp_aluResult~10_combout  & ((Mux91) # ((!Mux191 & Mux92))))

	.dataa(Mux19),
	.datab(Mux91),
	.datac(\temp_aluResult~10_combout ),
	.datad(Mux9),
	.cin(gnd),
	.combout(\temp_aluResult~26_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~26 .lut_mask = 16'h0F04;
defparam \temp_aluResult~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N16
cycloneive_lcell_comb \temp_aluResult~27 (
// Equation(s):
// \temp_aluResult~27_combout  = (!ex_mem_flush3 & (!temp_ALUop_output_3 & Mux61))

	.dataa(gnd),
	.datab(ex_mem_flush3),
	.datac(temp_ALUop_output_3),
	.datad(Mux6),
	.cin(gnd),
	.combout(\temp_aluResult~27_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~27 .lut_mask = 16'h0300;
defparam \temp_aluResult~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N22
cycloneive_lcell_comb \temp_aluResult~28 (
// Equation(s):
// \temp_aluResult~28_combout  = (!temp_ALUop_output_3 & (Mux71 & !ex_mem_flush3))

	.dataa(temp_ALUop_output_3),
	.datab(gnd),
	.datac(Mux7),
	.datad(ex_mem_flush3),
	.cin(gnd),
	.combout(\temp_aluResult~28_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~28 .lut_mask = 16'h0050;
defparam \temp_aluResult~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N12
cycloneive_lcell_comb \temp_aluResult~29 (
// Equation(s):
// \temp_aluResult~29_combout  = (!ex_mem_flush3 & (Mux51 & !temp_ALUop_output_3))

	.dataa(ex_mem_flush3),
	.datab(gnd),
	.datac(Mux5),
	.datad(temp_ALUop_output_3),
	.cin(gnd),
	.combout(\temp_aluResult~29_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~29 .lut_mask = 16'h0050;
defparam \temp_aluResult~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N8
cycloneive_lcell_comb \temp_aluResult~30 (
// Equation(s):
// \temp_aluResult~30_combout  = (!ex_mem_flush3 & (!temp_ALUop_output_3 & Mux41))

	.dataa(gnd),
	.datab(ex_mem_flush3),
	.datac(temp_ALUop_output_3),
	.datad(Mux4),
	.cin(gnd),
	.combout(\temp_aluResult~30_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~30 .lut_mask = 16'h0300;
defparam \temp_aluResult~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N18
cycloneive_lcell_comb \temp_aluResult~31 (
// Equation(s):
// \temp_aluResult~31_combout  = (!temp_ALUop_output_3 & (Mux210 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(temp_ALUop_output_3),
	.datac(Mux2),
	.datad(ex_mem_flush3),
	.cin(gnd),
	.combout(\temp_aluResult~31_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~31 .lut_mask = 16'h0030;
defparam \temp_aluResult~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N6
cycloneive_lcell_comb \temp_aluResult~32 (
// Equation(s):
// \temp_aluResult~32_combout  = (!\temp_aluResult~10_combout  & Mux32)

	.dataa(gnd),
	.datab(gnd),
	.datac(\temp_aluResult~10_combout ),
	.datad(Mux3),
	.cin(gnd),
	.combout(\temp_aluResult~32_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~32 .lut_mask = 16'h0F00;
defparam \temp_aluResult~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N6
cycloneive_lcell_comb \temp_aluResult~33 (
// Equation(s):
// \temp_aluResult~33_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux01)) # (!Mux191 & ((Mux02)))))

	.dataa(Mux0),
	.datab(\temp_aluResult~10_combout ),
	.datac(Mux19),
	.datad(Mux01),
	.cin(gnd),
	.combout(\temp_aluResult~33_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~33 .lut_mask = 16'h2320;
defparam \temp_aluResult~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N10
cycloneive_lcell_comb \temp_aluResult~34 (
// Equation(s):
// \temp_aluResult~34_combout  = (!\temp_aluResult~10_combout  & ((Mux191 & (Mux110)) # (!Mux191 & ((Mux113)))))

	.dataa(Mux1),
	.datab(Mux19),
	.datac(\temp_aluResult~10_combout ),
	.datad(Mux110),
	.cin(gnd),
	.combout(\temp_aluResult~34_combout ),
	.cout());
// synopsys translate_off
defparam \temp_aluResult~34 .lut_mask = 16'h0B08;
defparam \temp_aluResult~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N12
cycloneive_lcell_comb \temp_halt_out~0 (
// Equation(s):
// \temp_halt_out~0_combout  = (temp_halt_out_output1 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(temp_halt_out_output),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_halt_out~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_halt_out~0 .lut_mask = 16'h02AA;
defparam \temp_halt_out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N0
cycloneive_lcell_comb \temp_rdat2~60 (
// Equation(s):
// \temp_rdat2~60_combout  = (!ex_mem_flush3 & ((alu_b_mux_output_0) # (alu_b_mux_output_01)))

	.dataa(alu_b_mux_output_0),
	.datab(gnd),
	.datac(ex_mem_flush3),
	.datad(alu_b_mux_output_01),
	.cin(gnd),
	.combout(\temp_rdat2~60_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~60 .lut_mask = 16'h0F0A;
defparam \temp_rdat2~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N24
cycloneive_lcell_comb \temp_regwrite~0 (
// Equation(s):
// \temp_regwrite~0_combout  = (temp_regwrite_output1 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(temp_regwrite_output),
	.cin(gnd),
	.combout(\temp_regwrite~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_regwrite~0 .lut_mask = 16'h1F00;
defparam \temp_regwrite~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N6
cycloneive_lcell_comb \temp_memtoreg~0 (
// Equation(s):
// \temp_memtoreg~0_combout  = (temp_memtoreg_output_0 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(temp_memtoreg_output_0),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_memtoreg~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_memtoreg~0 .lut_mask = 16'h02AA;
defparam \temp_memtoreg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N6
cycloneive_lcell_comb \temp_memtoreg~1 (
// Equation(s):
// \temp_memtoreg~1_combout  = (temp_memtoreg_output_1 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(temp_memtoreg_output_1),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush2),
	.cin(gnd),
	.combout(\temp_memtoreg~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_memtoreg~1 .lut_mask = 16'h0A2A;
defparam \temp_memtoreg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N6
cycloneive_lcell_comb \temp_iMemLoad~0 (
// Equation(s):
// \temp_iMemLoad~0_combout  = (temp_imemload_output_0 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(temp_imemload_output_0),
	.cin(gnd),
	.combout(\temp_iMemLoad~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~0 .lut_mask = 16'h1F00;
defparam \temp_iMemLoad~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N20
cycloneive_lcell_comb \temp_iMemLoad~1 (
// Equation(s):
// \temp_iMemLoad~1_combout  = (temp_imemload_output_15 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(temp_imemload_output_15),
	.cin(gnd),
	.combout(\temp_iMemLoad~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~1 .lut_mask = 16'h3700;
defparam \temp_iMemLoad~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N22
cycloneive_lcell_comb \temp_iMemLoad~2 (
// Equation(s):
// \temp_iMemLoad~2_combout  = (temp_imemload_output_14 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(temp_imemload_output_14),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_iMemLoad~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~2 .lut_mask = 16'h222A;
defparam \temp_iMemLoad~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N4
cycloneive_lcell_comb \temp_iMemLoad~3 (
// Equation(s):
// \temp_iMemLoad~3_combout  = (temp_imemload_output_13 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(temp_imemload_output_13),
	.cin(gnd),
	.combout(\temp_iMemLoad~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~3 .lut_mask = 16'h1F00;
defparam \temp_iMemLoad~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N4
cycloneive_lcell_comb \temp_iMemLoad~4 (
// Equation(s):
// \temp_iMemLoad~4_combout  = (temp_imemload_output_10 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(temp_imemload_output_10),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_iMemLoad~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~4 .lut_mask = 16'h222A;
defparam \temp_iMemLoad~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N18
cycloneive_lcell_comb \temp_iMemLoad~5 (
// Equation(s):
// \temp_iMemLoad~5_combout  = (temp_imemload_output_9 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(temp_imemload_output_9),
	.cin(gnd),
	.combout(\temp_iMemLoad~5_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~5 .lut_mask = 16'h1F00;
defparam \temp_iMemLoad~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N4
cycloneive_lcell_comb \temp_iMemLoad~6 (
// Equation(s):
// \temp_iMemLoad~6_combout  = (temp_imemload_output_12 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(temp_imemload_output_12),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_iMemLoad~6_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~6 .lut_mask = 16'h10F0;
defparam \temp_iMemLoad~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N30
cycloneive_lcell_comb \temp_iMemLoad~7 (
// Equation(s):
// \temp_iMemLoad~7_combout  = (temp_imemload_output_11 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(temp_imemload_output_11),
	.cin(gnd),
	.combout(\temp_iMemLoad~7_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~7 .lut_mask = 16'h1F00;
defparam \temp_iMemLoad~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N16
cycloneive_lcell_comb \temp_iMemLoad~8 (
// Equation(s):
// \temp_iMemLoad~8_combout  = (temp_imemload_output_1 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(temp_imemload_output_1),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_iMemLoad~8_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~8 .lut_mask = 16'h10F0;
defparam \temp_iMemLoad~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N26
cycloneive_lcell_comb \temp_iMemLoad~9 (
// Equation(s):
// \temp_iMemLoad~9_combout  = (temp_imemload_output_4 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush),
	.datac(temp_imemload_output_4),
	.datad(ex_mem_flush2),
	.cin(gnd),
	.combout(\temp_iMemLoad~9_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~9 .lut_mask = 16'h3070;
defparam \temp_iMemLoad~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N30
cycloneive_lcell_comb \temp_iMemLoad~10 (
// Equation(s):
// \temp_iMemLoad~10_combout  = (temp_imemload_output_3 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(temp_imemload_output_3),
	.cin(gnd),
	.combout(\temp_iMemLoad~10_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~10 .lut_mask = 16'h3700;
defparam \temp_iMemLoad~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N16
cycloneive_lcell_comb \temp_iMemLoad~11 (
// Equation(s):
// \temp_iMemLoad~11_combout  = (temp_imemload_output_2 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(temp_imemload_output_2),
	.cin(gnd),
	.combout(\temp_iMemLoad~11_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~11 .lut_mask = 16'h3700;
defparam \temp_iMemLoad~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N4
cycloneive_lcell_comb \temp_iMemLoad~12 (
// Equation(s):
// \temp_iMemLoad~12_combout  = (temp_imemload_output_8 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(temp_imemload_output_8),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_iMemLoad~12_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~12 .lut_mask = 16'h10F0;
defparam \temp_iMemLoad~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N18
cycloneive_lcell_comb \temp_iMemLoad~13 (
// Equation(s):
// \temp_iMemLoad~13_combout  = (temp_imemload_output_7 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(temp_imemload_output_7),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_iMemLoad~13_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~13 .lut_mask = 16'h3070;
defparam \temp_iMemLoad~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N24
cycloneive_lcell_comb \temp_iMemLoad~14 (
// Equation(s):
// \temp_iMemLoad~14_combout  = (temp_imemload_output_6 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(temp_imemload_output_6),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_iMemLoad~14_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~14 .lut_mask = 16'h02AA;
defparam \temp_iMemLoad~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N22
cycloneive_lcell_comb \temp_iMemLoad~15 (
// Equation(s):
// \temp_iMemLoad~15_combout  = (temp_imemload_output_5 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(temp_imemload_output_5),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_iMemLoad~15_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~15 .lut_mask = 16'h444C;
defparam \temp_iMemLoad~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N6
cycloneive_lcell_comb \temp_iMemLoad~16 (
// Equation(s):
// \temp_iMemLoad~16_combout  = (temp_imemload_output_311 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(temp_imemload_output_31),
	.cin(gnd),
	.combout(\temp_iMemLoad~16_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~16 .lut_mask = 16'h3700;
defparam \temp_iMemLoad~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N28
cycloneive_lcell_comb \temp_iMemLoad~17 (
// Equation(s):
// \temp_iMemLoad~17_combout  = (temp_imemload_output_301 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(temp_imemload_output_30),
	.cin(gnd),
	.combout(\temp_iMemLoad~17_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~17 .lut_mask = 16'h3700;
defparam \temp_iMemLoad~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N24
cycloneive_lcell_comb \temp_iMemLoad~18 (
// Equation(s):
// \temp_iMemLoad~18_combout  = (temp_imemload_output_291 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(temp_imemload_output_29),
	.cin(gnd),
	.combout(\temp_iMemLoad~18_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~18 .lut_mask = 16'h3700;
defparam \temp_iMemLoad~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N0
cycloneive_lcell_comb \temp_iMemLoad~19 (
// Equation(s):
// \temp_iMemLoad~19_combout  = (temp_imemload_output_271 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(temp_imemload_output_27),
	.cin(gnd),
	.combout(\temp_iMemLoad~19_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~19 .lut_mask = 16'h3700;
defparam \temp_iMemLoad~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N18
cycloneive_lcell_comb \temp_iMemLoad~20 (
// Equation(s):
// \temp_iMemLoad~20_combout  = (temp_imemload_output_261 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(temp_imemload_output_26),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush1),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_iMemLoad~20_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~20 .lut_mask = 16'h02AA;
defparam \temp_iMemLoad~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N28
cycloneive_lcell_comb \temp_iMemLoad~21 (
// Equation(s):
// \temp_iMemLoad~21_combout  = (temp_imemload_output_281 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(temp_imemload_output_28),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_iMemLoad~21_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~21 .lut_mask = 16'h10F0;
defparam \temp_iMemLoad~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N2
cycloneive_lcell_comb \temp_branchSelect~0 (
// Equation(s):
// \temp_branchSelect~0_combout  = (temp_branch_output2 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(temp_branch_output),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_branchSelect~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_branchSelect~0 .lut_mask = 16'h0C4C;
defparam \temp_branchSelect~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N30
cycloneive_lcell_comb \temp_rdat1~63 (
// Equation(s):
// \temp_rdat1~63_combout  = (alu_a_mux_output_1 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush1),
	.datad(alu_a_mux_output_1),
	.cin(gnd),
	.combout(\temp_rdat1~63_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~63 .lut_mask = 16'h5700;
defparam \temp_rdat1~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N14
cycloneive_lcell_comb \temp_npc~0 (
// Equation(s):
// \temp_npc~0_combout  = (temp_NPC_output_1 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(temp_NPC_output_1),
	.cin(gnd),
	.combout(\temp_npc~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~0 .lut_mask = 16'h3700;
defparam \temp_npc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N0
cycloneive_lcell_comb \temp_pcselect~0 (
// Equation(s):
// \temp_pcselect~0_combout  = (temp_pcselect_output_1 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(temp_pcselect_output_1),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_pcselect~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_pcselect~0 .lut_mask = 16'h0C4C;
defparam \temp_pcselect~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N16
cycloneive_lcell_comb \temp_pcselect~1 (
// Equation(s):
// \temp_pcselect~1_combout  = (temp_pcselect_output_0 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush1),
	.datad(temp_pcselect_output_0),
	.cin(gnd),
	.combout(\temp_pcselect~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_pcselect~1 .lut_mask = 16'h5700;
defparam \temp_pcselect~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N8
cycloneive_lcell_comb \temp_rdat1~64 (
// Equation(s):
// \temp_rdat1~64_combout  = (alu_a_mux_output_0 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(alu_a_mux_output_0),
	.cin(gnd),
	.combout(\temp_rdat1~64_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~64 .lut_mask = 16'h3700;
defparam \temp_rdat1~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N28
cycloneive_lcell_comb \temp_npc~1 (
// Equation(s):
// \temp_npc~1_combout  = (temp_NPC_output_0 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(temp_NPC_output_0),
	.cin(gnd),
	.combout(\temp_npc~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~1 .lut_mask = 16'h3700;
defparam \temp_npc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N18
cycloneive_lcell_comb \temp_npc~2 (
// Equation(s):
// \temp_npc~2_combout  = (temp_NPC_output_2 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(temp_NPC_output_2),
	.cin(gnd),
	.combout(\temp_npc~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~2 .lut_mask = 16'h3700;
defparam \temp_npc~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N24
cycloneive_lcell_comb \temp_rdat1~65 (
// Equation(s):
// \temp_rdat1~65_combout  = (alu_a_mux_output_2 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(alu_a_mux_output_2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~65_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~65 .lut_mask = 16'h3070;
defparam \temp_rdat1~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N10
cycloneive_lcell_comb \temp_npc~3 (
// Equation(s):
// \temp_npc~3_combout  = (temp_NPC_output_3 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush1),
	.datad(temp_NPC_output_3),
	.cin(gnd),
	.combout(\temp_npc~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~3 .lut_mask = 16'h5700;
defparam \temp_npc~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N22
cycloneive_lcell_comb \temp_rdat1~62 (
// Equation(s):
// \temp_rdat1~62_combout  = (!ex_mem_flush3 & ((alu_a_mux_output_32) # (alu_a_mux_output_3)))

	.dataa(ex_mem_flush3),
	.datab(gnd),
	.datac(alu_a_mux_output_32),
	.datad(alu_a_mux_output_3),
	.cin(gnd),
	.combout(\temp_rdat1~62_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~62 .lut_mask = 16'h5550;
defparam \temp_rdat1~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N14
cycloneive_lcell_comb \temp_npc~4 (
// Equation(s):
// \temp_npc~4_combout  = (temp_NPC_output_5 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(temp_NPC_output_5),
	.cin(gnd),
	.combout(\temp_npc~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~4 .lut_mask = 16'h3700;
defparam \temp_npc~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N0
cycloneive_lcell_comb \temp_npc~5 (
// Equation(s):
// \temp_npc~5_combout  = (temp_NPC_output_4 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(temp_NPC_output_4),
	.cin(gnd),
	.combout(\temp_npc~5_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~5 .lut_mask = 16'h3700;
defparam \temp_npc~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N28
cycloneive_lcell_comb \temp_rdat1~66 (
// Equation(s):
// \temp_rdat1~66_combout  = (alu_a_mux_output_5 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(alu_a_mux_output_5),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~66_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~66 .lut_mask = 16'h5070;
defparam \temp_rdat1~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N10
cycloneive_lcell_comb \temp_rdat1~67 (
// Equation(s):
// \temp_rdat1~67_combout  = (alu_a_mux_output_4 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(alu_a_mux_output_4),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~67_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~67 .lut_mask = 16'h3070;
defparam \temp_rdat1~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N2
cycloneive_lcell_comb \temp_npc~6 (
// Equation(s):
// \temp_npc~6_combout  = (temp_NPC_output_7 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(temp_NPC_output_7),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_npc~6_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~6 .lut_mask = 16'h0A2A;
defparam \temp_npc~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N20
cycloneive_lcell_comb \temp_npc~7 (
// Equation(s):
// \temp_npc~7_combout  = (temp_NPC_output_6 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush1),
	.datad(temp_NPC_output_6),
	.cin(gnd),
	.combout(\temp_npc~7_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~7 .lut_mask = 16'h5700;
defparam \temp_npc~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N24
cycloneive_lcell_comb \temp_rdat1~68 (
// Equation(s):
// \temp_rdat1~68_combout  = (alu_a_mux_output_7 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(alu_a_mux_output_7),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~68_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~68 .lut_mask = 16'h0A2A;
defparam \temp_rdat1~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N2
cycloneive_lcell_comb \temp_rdat1~69 (
// Equation(s):
// \temp_rdat1~69_combout  = (alu_a_mux_output_6 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(alu_a_mux_output_6),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~69_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~69 .lut_mask = 16'h3070;
defparam \temp_rdat1~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y45_N0
cycloneive_lcell_comb \temp_rdat1[6]~feeder (
// Equation(s):
// \temp_rdat1[6]~feeder_combout  = \temp_rdat1~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\temp_rdat1~69_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_rdat1[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1[6]~feeder .lut_mask = 16'hF0F0;
defparam \temp_rdat1[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N8
cycloneive_lcell_comb \temp_npc~8 (
// Equation(s):
// \temp_npc~8_combout  = (temp_NPC_output_9 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(temp_NPC_output_9),
	.cin(gnd),
	.combout(\temp_npc~8_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~8 .lut_mask = 16'h3700;
defparam \temp_npc~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N28
cycloneive_lcell_comb \temp_npc~9 (
// Equation(s):
// \temp_npc~9_combout  = (temp_NPC_output_8 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(temp_NPC_output_8),
	.cin(gnd),
	.combout(\temp_npc~9_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~9 .lut_mask = 16'h1F00;
defparam \temp_npc~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N6
cycloneive_lcell_comb \temp_rdat1~70 (
// Equation(s):
// \temp_rdat1~70_combout  = (alu_a_mux_output_9 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(alu_a_mux_output_9),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_rdat1~70_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~70 .lut_mask = 16'h04CC;
defparam \temp_rdat1~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N6
cycloneive_lcell_comb \temp_rdat1~71 (
// Equation(s):
// \temp_rdat1~71_combout  = (alu_a_mux_output_8 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(alu_a_mux_output_8),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~71_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~71 .lut_mask = 16'h3070;
defparam \temp_rdat1~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N18
cycloneive_lcell_comb \temp_npc~10 (
// Equation(s):
// \temp_npc~10_combout  = (temp_NPC_output_11 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(temp_NPC_output_11),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_npc~10_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~10 .lut_mask = 16'h444C;
defparam \temp_npc~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N18
cycloneive_lcell_comb \temp_npc~11 (
// Equation(s):
// \temp_npc~11_combout  = (temp_NPC_output_10 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(temp_NPC_output_10),
	.cin(gnd),
	.combout(\temp_npc~11_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~11 .lut_mask = 16'h1F00;
defparam \temp_npc~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N0
cycloneive_lcell_comb \temp_rdat1~72 (
// Equation(s):
// \temp_rdat1~72_combout  = (alu_a_mux_output_11 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(alu_a_mux_output_11),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_rdat1~72_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~72 .lut_mask = 16'h10F0;
defparam \temp_rdat1~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N16
cycloneive_lcell_comb \temp_rdat1~73 (
// Equation(s):
// \temp_rdat1~73_combout  = (alu_a_mux_output_10 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(alu_a_mux_output_10),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~73_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~73 .lut_mask = 16'h0C4C;
defparam \temp_rdat1~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N0
cycloneive_lcell_comb \temp_npc~12 (
// Equation(s):
// \temp_npc~12_combout  = (temp_NPC_output_13 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(temp_NPC_output_13),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_npc~12_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~12 .lut_mask = 16'h10F0;
defparam \temp_npc~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N8
cycloneive_lcell_comb \temp_npc~13 (
// Equation(s):
// \temp_npc~13_combout  = (temp_NPC_output_12 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(temp_NPC_output_12),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_npc~13_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~13 .lut_mask = 16'h10F0;
defparam \temp_npc~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N16
cycloneive_lcell_comb \temp_rdat1~74 (
// Equation(s):
// \temp_rdat1~74_combout  = (alu_a_mux_output_13 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(alu_a_mux_output_13),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_rdat1~74_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~74 .lut_mask = 16'h02AA;
defparam \temp_rdat1~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N26
cycloneive_lcell_comb \temp_rdat1~75 (
// Equation(s):
// \temp_rdat1~75_combout  = (alu_a_mux_output_12 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(alu_a_mux_output_12),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~75_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~75 .lut_mask = 16'h0C4C;
defparam \temp_rdat1~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N24
cycloneive_lcell_comb \temp_npc~14 (
// Equation(s):
// \temp_npc~14_combout  = (temp_NPC_output_15 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(temp_NPC_output_15),
	.cin(gnd),
	.combout(\temp_npc~14_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~14 .lut_mask = 16'h1F00;
defparam \temp_npc~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N22
cycloneive_lcell_comb \temp_npc~15 (
// Equation(s):
// \temp_npc~15_combout  = (temp_NPC_output_14 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(temp_NPC_output_14),
	.cin(gnd),
	.combout(\temp_npc~15_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~15 .lut_mask = 16'h1F00;
defparam \temp_npc~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N12
cycloneive_lcell_comb \temp_rdat1~76 (
// Equation(s):
// \temp_rdat1~76_combout  = (alu_a_mux_output_15 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(alu_a_mux_output_15),
	.cin(gnd),
	.combout(\temp_rdat1~76_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~76 .lut_mask = 16'h5700;
defparam \temp_rdat1~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N2
cycloneive_lcell_comb \temp_rdat1~77 (
// Equation(s):
// \temp_rdat1~77_combout  = (alu_a_mux_output_14 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(alu_a_mux_output_14),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~77_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~77 .lut_mask = 16'h3070;
defparam \temp_rdat1~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N20
cycloneive_lcell_comb \temp_npc~16 (
// Equation(s):
// \temp_npc~16_combout  = (temp_NPC_output_17 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(temp_NPC_output_17),
	.cin(gnd),
	.combout(\temp_npc~16_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~16 .lut_mask = 16'h5700;
defparam \temp_npc~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N2
cycloneive_lcell_comb \temp_npc~17 (
// Equation(s):
// \temp_npc~17_combout  = (temp_NPC_output_16 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(temp_NPC_output_16),
	.cin(gnd),
	.combout(\temp_npc~17_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~17 .lut_mask = 16'h1F00;
defparam \temp_npc~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N8
cycloneive_lcell_comb \temp_rdat1~78 (
// Equation(s):
// \temp_rdat1~78_combout  = (alu_a_mux_output_17 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush1),
	.datad(alu_a_mux_output_17),
	.cin(gnd),
	.combout(\temp_rdat1~78_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~78 .lut_mask = 16'h5700;
defparam \temp_rdat1~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N8
cycloneive_lcell_comb \temp_rdat1~79 (
// Equation(s):
// \temp_rdat1~79_combout  = (alu_a_mux_output_16 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(alu_a_mux_output_16),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_rdat1~79_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~79 .lut_mask = 16'h04CC;
defparam \temp_rdat1~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N2
cycloneive_lcell_comb \temp_signZero~0 (
// Equation(s):
// \temp_signZero~0_combout  = (temp_signzerovalue_output_16 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(temp_signzerovalue_output_16),
	.cin(gnd),
	.combout(\temp_signZero~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_signZero~0 .lut_mask = 16'h1F00;
defparam \temp_signZero~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N28
cycloneive_lcell_comb \temp_npc~18 (
// Equation(s):
// \temp_npc~18_combout  = (temp_NPC_output_19 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(temp_NPC_output_19),
	.cin(gnd),
	.combout(\temp_npc~18_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~18 .lut_mask = 16'h3700;
defparam \temp_npc~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N4
cycloneive_lcell_comb \temp_npc~19 (
// Equation(s):
// \temp_npc~19_combout  = (temp_NPC_output_18 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush1),
	.datad(temp_NPC_output_18),
	.cin(gnd),
	.combout(\temp_npc~19_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~19 .lut_mask = 16'h5700;
defparam \temp_npc~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N0
cycloneive_lcell_comb \temp_rdat1~80 (
// Equation(s):
// \temp_rdat1~80_combout  = (alu_a_mux_output_19 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(alu_a_mux_output_19),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~80_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~80 .lut_mask = 16'h3070;
defparam \temp_rdat1~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N0
cycloneive_lcell_comb \temp_iMemLoad~22 (
// Equation(s):
// \temp_iMemLoad~22_combout  = (temp_imemload_output_17 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\temp_iMemLoad~22_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~22 .lut_mask = 16'h3700;
defparam \temp_iMemLoad~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N14
cycloneive_lcell_comb \temp_rdat1~81 (
// Equation(s):
// \temp_rdat1~81_combout  = (alu_a_mux_output_18 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(alu_a_mux_output_18),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_rdat1~81_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~81 .lut_mask = 16'h04CC;
defparam \temp_rdat1~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N14
cycloneive_lcell_comb \temp_iMemLoad~23 (
// Equation(s):
// \temp_iMemLoad~23_combout  = (temp_imemload_output_16 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(temp_imemload_output_16),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_iMemLoad~23_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~23 .lut_mask = 16'h0C4C;
defparam \temp_iMemLoad~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N6
cycloneive_lcell_comb \temp_npc~20 (
// Equation(s):
// \temp_npc~20_combout  = (temp_NPC_output_20 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(temp_NPC_output_20),
	.cin(gnd),
	.combout(\temp_npc~20_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~20 .lut_mask = 16'h5700;
defparam \temp_npc~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N2
cycloneive_lcell_comb \temp_rdat1~82 (
// Equation(s):
// \temp_rdat1~82_combout  = (alu_a_mux_output_20 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(alu_a_mux_output_20),
	.cin(gnd),
	.combout(\temp_rdat1~82_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~82 .lut_mask = 16'h1F00;
defparam \temp_rdat1~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N0
cycloneive_lcell_comb \temp_iMemLoad~24 (
// Equation(s):
// \temp_iMemLoad~24_combout  = (temp_imemload_output_18 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(temp_imemload_output_18),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_iMemLoad~24_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~24 .lut_mask = 16'h02AA;
defparam \temp_iMemLoad~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N12
cycloneive_lcell_comb \temp_npc~21 (
// Equation(s):
// \temp_npc~21_combout  = (temp_NPC_output_21 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(temp_NPC_output_21),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_npc~21_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~21 .lut_mask = 16'h02AA;
defparam \temp_npc~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N8
cycloneive_lcell_comb \temp_rdat1~83 (
// Equation(s):
// \temp_rdat1~83_combout  = (alu_a_mux_output_21 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(alu_a_mux_output_21),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~83_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~83 .lut_mask = 16'h3070;
defparam \temp_rdat1~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N4
cycloneive_lcell_comb \temp_iMemLoad~25 (
// Equation(s):
// \temp_iMemLoad~25_combout  = (temp_imemload_output_19 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(temp_imemload_output_19),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_iMemLoad~25_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~25 .lut_mask = 16'h222A;
defparam \temp_iMemLoad~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N2
cycloneive_lcell_comb \temp_npc~22 (
// Equation(s):
// \temp_npc~22_combout  = (temp_NPC_output_23 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(temp_NPC_output_23),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(ex_mem_flush2),
	.cin(gnd),
	.combout(\temp_npc~22_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~22 .lut_mask = 16'h222A;
defparam \temp_npc~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y44_N30
cycloneive_lcell_comb \temp_npc~23 (
// Equation(s):
// \temp_npc~23_combout  = (temp_NPC_output_22 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(temp_NPC_output_22),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_npc~23_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~23 .lut_mask = 16'h02AA;
defparam \temp_npc~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N18
cycloneive_lcell_comb \temp_rdat1~84 (
// Equation(s):
// \temp_rdat1~84_combout  = (alu_a_mux_output_23 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(alu_a_mux_output_23),
	.cin(gnd),
	.combout(\temp_rdat1~84_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~84 .lut_mask = 16'h3700;
defparam \temp_rdat1~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N2
cycloneive_lcell_comb \temp_iMemLoad~26 (
// Equation(s):
// \temp_iMemLoad~26_combout  = (temp_imemload_output_21 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(temp_imemload_output_21),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_iMemLoad~26_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~26 .lut_mask = 16'h3070;
defparam \temp_iMemLoad~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N2
cycloneive_lcell_comb \temp_rdat1~85 (
// Equation(s):
// \temp_rdat1~85_combout  = (alu_a_mux_output_22 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(alu_a_mux_output_22),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~85_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~85 .lut_mask = 16'h5070;
defparam \temp_rdat1~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N10
cycloneive_lcell_comb \temp_iMemLoad~27 (
// Equation(s):
// \temp_iMemLoad~27_combout  = (temp_imemload_output_20 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(temp_imemload_output_20),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_iMemLoad~27_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~27 .lut_mask = 16'h5070;
defparam \temp_iMemLoad~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N12
cycloneive_lcell_comb \temp_npc~24 (
// Equation(s):
// \temp_npc~24_combout  = (temp_NPC_output_25 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(temp_NPC_output_25),
	.cin(gnd),
	.combout(\temp_npc~24_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~24 .lut_mask = 16'h3700;
defparam \temp_npc~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N10
cycloneive_lcell_comb \temp_npc~25 (
// Equation(s):
// \temp_npc~25_combout  = (temp_NPC_output_24 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(temp_NPC_output_24),
	.cin(gnd),
	.combout(\temp_npc~25_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~25 .lut_mask = 16'h3700;
defparam \temp_npc~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N0
cycloneive_lcell_comb \temp_rdat1~86 (
// Equation(s):
// \temp_rdat1~86_combout  = (alu_a_mux_output_25 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(alu_a_mux_output_25),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~86_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~86 .lut_mask = 16'h0C4C;
defparam \temp_rdat1~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N14
cycloneive_lcell_comb \temp_iMemLoad~28 (
// Equation(s):
// \temp_iMemLoad~28_combout  = (temp_imemload_output_23 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(temp_imemload_output_23),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_iMemLoad~28_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~28 .lut_mask = 16'h0C4C;
defparam \temp_iMemLoad~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N6
cycloneive_lcell_comb \temp_rdat1~87 (
// Equation(s):
// \temp_rdat1~87_combout  = (alu_a_mux_output_24 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(alu_a_mux_output_24),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush1),
	.datad(ex_mem_flush2),
	.cin(gnd),
	.combout(\temp_rdat1~87_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~87 .lut_mask = 16'h222A;
defparam \temp_rdat1~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N30
cycloneive_lcell_comb \temp_iMemLoad~29 (
// Equation(s):
// \temp_iMemLoad~29_combout  = (temp_imemload_output_22 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(temp_imemload_output_22),
	.datac(ex_mem_flush1),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_iMemLoad~29_combout ),
	.cout());
// synopsys translate_off
defparam \temp_iMemLoad~29 .lut_mask = 16'h04CC;
defparam \temp_iMemLoad~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N2
cycloneive_lcell_comb \temp_npc~26 (
// Equation(s):
// \temp_npc~26_combout  = (temp_NPC_output_26 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(temp_NPC_output_26),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_npc~26_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~26 .lut_mask = 16'h444C;
defparam \temp_npc~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N8
cycloneive_lcell_comb \temp_rdat1~88 (
// Equation(s):
// \temp_rdat1~88_combout  = (alu_a_mux_output_26 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(alu_a_mux_output_26),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~88_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~88 .lut_mask = 16'h0C4C;
defparam \temp_rdat1~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N4
cycloneive_lcell_comb \temp_npc~27 (
// Equation(s):
// \temp_npc~27_combout  = (temp_NPC_output_27 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(temp_NPC_output_27),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_npc~27_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~27 .lut_mask = 16'h444C;
defparam \temp_npc~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N18
cycloneive_lcell_comb \temp_rdat1~89 (
// Equation(s):
// \temp_rdat1~89_combout  = (alu_a_mux_output_27 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(alu_a_mux_output_27),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_rdat1~89_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~89 .lut_mask = 16'h10F0;
defparam \temp_rdat1~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N18
cycloneive_lcell_comb \temp_npc~28 (
// Equation(s):
// \temp_npc~28_combout  = (temp_NPC_output_29 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(temp_NPC_output_29),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_npc~28_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~28 .lut_mask = 16'h444C;
defparam \temp_npc~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N10
cycloneive_lcell_comb \temp_npc~29 (
// Equation(s):
// \temp_npc~29_combout  = (temp_NPC_output_28 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(temp_NPC_output_28),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_npc~29_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~29 .lut_mask = 16'h444C;
defparam \temp_npc~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N22
cycloneive_lcell_comb \temp_rdat1~90 (
// Equation(s):
// \temp_rdat1~90_combout  = (alu_a_mux_output_29 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(alu_a_mux_output_29),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~90_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~90 .lut_mask = 16'h5070;
defparam \temp_rdat1~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N12
cycloneive_lcell_comb \temp_rdat1~91 (
// Equation(s):
// \temp_rdat1~91_combout  = (alu_a_mux_output_28 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(alu_a_mux_output_28),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat1~91_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~91 .lut_mask = 16'h444C;
defparam \temp_rdat1~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N18
cycloneive_lcell_comb \temp_rdat1~92 (
// Equation(s):
// \temp_rdat1~92_combout  = (alu_a_mux_output_311 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(alu_a_mux_output_31),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_rdat1~92_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~92 .lut_mask = 16'h02AA;
defparam \temp_rdat1~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N30
cycloneive_lcell_comb \temp_npc~30 (
// Equation(s):
// \temp_npc~30_combout  = (temp_NPC_output_31 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(temp_NPC_output_31),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_npc~30_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~30 .lut_mask = 16'h10F0;
defparam \temp_npc~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N12
cycloneive_lcell_comb \temp_npc~31 (
// Equation(s):
// \temp_npc~31_combout  = (temp_NPC_output_30 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(temp_NPC_output_30),
	.cin(gnd),
	.combout(\temp_npc~31_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc~31 .lut_mask = 16'h1F00;
defparam \temp_npc~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N12
cycloneive_lcell_comb \temp_rdat1~93 (
// Equation(s):
// \temp_rdat1~93_combout  = (alu_a_mux_output_30 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush1),
	.datad(alu_a_mux_output_30),
	.cin(gnd),
	.combout(\temp_rdat1~93_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat1~93 .lut_mask = 16'h5700;
defparam \temp_rdat1~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N6
cycloneive_lcell_comb \temp_rdat2~61 (
// Equation(s):
// \temp_rdat2~61_combout  = (!ex_mem_flush3 & ((alu_b_mux_output_11) # (alu_b_mux_output_1)))

	.dataa(gnd),
	.datab(alu_b_mux_output_11),
	.datac(ex_mem_flush3),
	.datad(alu_b_mux_output_1),
	.cin(gnd),
	.combout(\temp_rdat2~61_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~61 .lut_mask = 16'h0F0C;
defparam \temp_rdat2~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N28
cycloneive_lcell_comb \temp_rdat2~62 (
// Equation(s):
// \temp_rdat2~62_combout  = (alu_b_mux_output_2 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(alu_b_mux_output_2),
	.cin(gnd),
	.combout(\temp_rdat2~62_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~62 .lut_mask = 16'h1F00;
defparam \temp_rdat2~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N4
cycloneive_lcell_comb \temp_rdat2~63 (
// Equation(s):
// \temp_rdat2~63_combout  = (alu_b_mux_output_3 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(alu_b_mux_output_3),
	.cin(gnd),
	.combout(\temp_rdat2~63_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~63 .lut_mask = 16'h5700;
defparam \temp_rdat2~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N16
cycloneive_lcell_comb \temp_rdat2~64 (
// Equation(s):
// \temp_rdat2~64_combout  = (alu_b_mux_output_4 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(alu_b_mux_output_4),
	.cin(gnd),
	.combout(\temp_rdat2~64_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~64 .lut_mask = 16'h1F00;
defparam \temp_rdat2~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N14
cycloneive_lcell_comb \temp_rdat2~65 (
// Equation(s):
// \temp_rdat2~65_combout  = (alu_b_mux_output_5 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(alu_b_mux_output_5),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat2~65_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~65 .lut_mask = 16'h444C;
defparam \temp_rdat2~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N30
cycloneive_lcell_comb \temp_rdat2~66 (
// Equation(s):
// \temp_rdat2~66_combout  = (alu_b_mux_output_6 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(alu_b_mux_output_6),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat2~66_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~66 .lut_mask = 16'h3070;
defparam \temp_rdat2~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N14
cycloneive_lcell_comb \temp_rdat2~67 (
// Equation(s):
// \temp_rdat2~67_combout  = (alu_b_mux_output_7 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(alu_b_mux_output_7),
	.cin(gnd),
	.combout(\temp_rdat2~67_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~67 .lut_mask = 16'h1F00;
defparam \temp_rdat2~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N10
cycloneive_lcell_comb \temp_rdat2~68 (
// Equation(s):
// \temp_rdat2~68_combout  = (alu_b_mux_output_8 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(alu_b_mux_output_8),
	.cin(gnd),
	.combout(\temp_rdat2~68_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~68 .lut_mask = 16'h1F00;
defparam \temp_rdat2~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N20
cycloneive_lcell_comb \temp_rdat2~69 (
// Equation(s):
// \temp_rdat2~69_combout  = (alu_b_mux_output_9 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(alu_b_mux_output_9),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush2),
	.cin(gnd),
	.combout(\temp_rdat2~69_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~69 .lut_mask = 16'h0A2A;
defparam \temp_rdat2~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N8
cycloneive_lcell_comb \temp_rdat2~70 (
// Equation(s):
// \temp_rdat2~70_combout  = (alu_b_mux_output_10 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(alu_b_mux_output_10),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush2),
	.cin(gnd),
	.combout(\temp_rdat2~70_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~70 .lut_mask = 16'h0C4C;
defparam \temp_rdat2~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N24
cycloneive_lcell_comb \temp_rdat2~71 (
// Equation(s):
// \temp_rdat2~71_combout  = (alu_b_mux_output_111 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(alu_b_mux_output_111),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat2~71_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~71 .lut_mask = 16'h3070;
defparam \temp_rdat2~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N2
cycloneive_lcell_comb \temp_rdat2~72 (
// Equation(s):
// \temp_rdat2~72_combout  = (alu_b_mux_output_12 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(alu_b_mux_output_12),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat2~72_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~72 .lut_mask = 16'h5070;
defparam \temp_rdat2~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N26
cycloneive_lcell_comb \temp_rdat2~73 (
// Equation(s):
// \temp_rdat2~73_combout  = (alu_b_mux_output_13 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(alu_b_mux_output_13),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat2~73_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~73 .lut_mask = 16'h444C;
defparam \temp_rdat2~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N20
cycloneive_lcell_comb \temp_rdat2~74 (
// Equation(s):
// \temp_rdat2~74_combout  = (alu_b_mux_output_14 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(alu_b_mux_output_14),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat2~74_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~74 .lut_mask = 16'h3070;
defparam \temp_rdat2~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N26
cycloneive_lcell_comb \temp_rdat2~75 (
// Equation(s):
// \temp_rdat2~75_combout  = (alu_b_mux_output_15 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(alu_b_mux_output_15),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush2),
	.cin(gnd),
	.combout(\temp_rdat2~75_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~75 .lut_mask = 16'h0A2A;
defparam \temp_rdat2~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N30
cycloneive_lcell_comb \temp_rdat2~76 (
// Equation(s):
// \temp_rdat2~76_combout  = (alu_b_mux_output_16 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(alu_b_mux_output_16),
	.cin(gnd),
	.combout(\temp_rdat2~76_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~76 .lut_mask = 16'h1F00;
defparam \temp_rdat2~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N18
cycloneive_lcell_comb \temp_rdat2~77 (
// Equation(s):
// \temp_rdat2~77_combout  = (alu_b_mux_output_17 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(alu_b_mux_output_17),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat2~77_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~77 .lut_mask = 16'h0A2A;
defparam \temp_rdat2~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N24
cycloneive_lcell_comb \temp_rdat2~78 (
// Equation(s):
// \temp_rdat2~78_combout  = (alu_b_mux_output_18 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(alu_b_mux_output_18),
	.cin(gnd),
	.combout(\temp_rdat2~78_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~78 .lut_mask = 16'h1F00;
defparam \temp_rdat2~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N30
cycloneive_lcell_comb \temp_rdat2~79 (
// Equation(s):
// \temp_rdat2~79_combout  = (alu_b_mux_output_19 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(alu_b_mux_output_19),
	.cin(gnd),
	.combout(\temp_rdat2~79_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~79 .lut_mask = 16'h1F00;
defparam \temp_rdat2~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N8
cycloneive_lcell_comb \temp_rdat2~80 (
// Equation(s):
// \temp_rdat2~80_combout  = (alu_b_mux_output_20 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(alu_b_mux_output_20),
	.cin(gnd),
	.combout(\temp_rdat2~80_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~80 .lut_mask = 16'h1F00;
defparam \temp_rdat2~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N26
cycloneive_lcell_comb \temp_rdat2~81 (
// Equation(s):
// \temp_rdat2~81_combout  = (alu_b_mux_output_21 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(alu_b_mux_output_21),
	.cin(gnd),
	.combout(\temp_rdat2~81_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~81 .lut_mask = 16'h1F00;
defparam \temp_rdat2~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N26
cycloneive_lcell_comb \temp_rdat2~82 (
// Equation(s):
// \temp_rdat2~82_combout  = (alu_b_mux_output_22 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush1),
	.datad(alu_b_mux_output_22),
	.cin(gnd),
	.combout(\temp_rdat2~82_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~82 .lut_mask = 16'h5700;
defparam \temp_rdat2~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N24
cycloneive_lcell_comb \temp_rdat2~83 (
// Equation(s):
// \temp_rdat2~83_combout  = (alu_b_mux_output_23 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(alu_b_mux_output_23),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_rdat2~83_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~83 .lut_mask = 16'h04CC;
defparam \temp_rdat2~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N24
cycloneive_lcell_comb \temp_rdat2~84 (
// Equation(s):
// \temp_rdat2~84_combout  = (alu_b_mux_output_24 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(alu_b_mux_output_24),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat2~84_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~84 .lut_mask = 16'h0A2A;
defparam \temp_rdat2~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N10
cycloneive_lcell_comb \temp_rdat2~85 (
// Equation(s):
// \temp_rdat2~85_combout  = (alu_b_mux_output_25 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(alu_b_mux_output_25),
	.cin(gnd),
	.combout(\temp_rdat2~85_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~85 .lut_mask = 16'h1F00;
defparam \temp_rdat2~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N22
cycloneive_lcell_comb \temp_rdat2~86 (
// Equation(s):
// \temp_rdat2~86_combout  = (alu_b_mux_output_26 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(alu_b_mux_output_26),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat2~86_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~86 .lut_mask = 16'h0C4C;
defparam \temp_rdat2~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N28
cycloneive_lcell_comb \temp_rdat2~87 (
// Equation(s):
// \temp_rdat2~87_combout  = (alu_b_mux_output_27 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush),
	.datac(alu_b_mux_output_27),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat2~87_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~87 .lut_mask = 16'h3070;
defparam \temp_rdat2~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N16
cycloneive_lcell_comb \temp_rdat2~88 (
// Equation(s):
// \temp_rdat2~88_combout  = (alu_b_mux_output_28 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(alu_b_mux_output_28),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_rdat2~88_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~88 .lut_mask = 16'h02AA;
defparam \temp_rdat2~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N14
cycloneive_lcell_comb \temp_rdat2~89 (
// Equation(s):
// \temp_rdat2~89_combout  = (alu_b_mux_output_29 & (((!ex_mem_flush1 & !ex_mem_flush2)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush1),
	.datab(alu_b_mux_output_29),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush2),
	.cin(gnd),
	.combout(\temp_rdat2~89_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~89 .lut_mask = 16'h0C4C;
defparam \temp_rdat2~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N18
cycloneive_lcell_comb \temp_rdat2~90 (
// Equation(s):
// \temp_rdat2~90_combout  = (alu_b_mux_output_30 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(ex_mem_flush2),
	.datab(ex_mem_flush1),
	.datac(ex_mem_flush),
	.datad(alu_b_mux_output_30),
	.cin(gnd),
	.combout(\temp_rdat2~90_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~90 .lut_mask = 16'h1F00;
defparam \temp_rdat2~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N6
cycloneive_lcell_comb \temp_rdat2~91 (
// Equation(s):
// \temp_rdat2~91_combout  = (alu_b_mux_output_31 & (((!ex_mem_flush2 & !ex_mem_flush1)) # (!ex_mem_flush)))

	.dataa(alu_b_mux_output_31),
	.datab(ex_mem_flush2),
	.datac(ex_mem_flush),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(\temp_rdat2~91_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat2~91 .lut_mask = 16'h0A2A;
defparam \temp_rdat2~91 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module extender (
	temp_imemload_output_31,
	temp_imemload_output_30,
	Equal3,
	temp_branch_output,
	temp_imemload_output_15,
	Equal31,
	extended_imm_16,
	temp_ALUsrc_output,
	WideOr5,
	extended_imm_161,
	devpor,
	devclrn,
	devoe);
input 	temp_imemload_output_31;
input 	temp_imemload_output_30;
input 	Equal3;
input 	temp_branch_output;
input 	temp_imemload_output_15;
input 	Equal31;
output 	extended_imm_16;
input 	temp_ALUsrc_output;
input 	WideOr5;
output 	extended_imm_161;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \extended_imm[16]~1_combout ;


// Location: LCCOMB_X65_Y37_N6
cycloneive_lcell_comb \extended_imm[16]~0 (
// Equation(s):
// extended_imm_16 = (!temp_imemload_output_30 & (((Equal32) # (!Equal3)) # (!temp_branch_output1)))

	.dataa(temp_branch_output),
	.datab(temp_imemload_output_30),
	.datac(Equal3),
	.datad(Equal31),
	.cin(gnd),
	.combout(extended_imm_16),
	.cout());
// synopsys translate_off
defparam \extended_imm[16]~0 .lut_mask = 16'h3313;
defparam \extended_imm[16]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N20
cycloneive_lcell_comb \extended_imm[16]~2 (
// Equation(s):
// extended_imm_161 = (\extended_imm[16]~1_combout  & extended_imm_16)

	.dataa(gnd),
	.datab(\extended_imm[16]~1_combout ),
	.datac(extended_imm_16),
	.datad(gnd),
	.cin(gnd),
	.combout(extended_imm_161),
	.cout());
// synopsys translate_off
defparam \extended_imm[16]~2 .lut_mask = 16'hC0C0;
defparam \extended_imm[16]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N4
cycloneive_lcell_comb \extended_imm[16]~1 (
// Equation(s):
// \extended_imm[16]~1_combout  = (temp_imemload_output_15 & ((temp_ALUsrc_output) # ((WideOr5 & !temp_imemload_output_31))))

	.dataa(WideOr5),
	.datab(temp_ALUsrc_output),
	.datac(temp_imemload_output_31),
	.datad(temp_imemload_output_15),
	.cin(gnd),
	.combout(\extended_imm[16]~1_combout ),
	.cout());
// synopsys translate_off
defparam \extended_imm[16]~1 .lut_mask = 16'hCE00;
defparam \extended_imm[16]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module forward (
	temp_branchDest_0,
	temp_branchDest_4,
	temp_branchDest_3,
	temp_branchDest_2,
	temp_branchDest_1,
	temp_regwrite,
	temp_imemload_output_17,
	temp_imemload_output_16,
	temp_imemload_output_18,
	temp_imemload_output_19,
	temp_imemload_output_20,
	temp_memtoreg_0,
	temp_memtoreg_1,
	always0,
	temp_regwrite1,
	always01,
	temp_branchDest_11,
	temp_branchDest_01,
	temp_branchDest_31,
	temp_branchDest_21,
	temp_branchDest_41,
	always02,
	always03,
	forwardb_1,
	temp_imemload_output_22,
	temp_imemload_output_21,
	temp_imemload_output_23,
	temp_imemload_output_24,
	temp_imemload_output_25,
	forwarda_1,
	always04,
	always05,
	always06,
	always07,
	devpor,
	devclrn,
	devoe);
input 	temp_branchDest_0;
input 	temp_branchDest_4;
input 	temp_branchDest_3;
input 	temp_branchDest_2;
input 	temp_branchDest_1;
input 	temp_regwrite;
input 	temp_imemload_output_17;
input 	temp_imemload_output_16;
input 	temp_imemload_output_18;
input 	temp_imemload_output_19;
input 	temp_imemload_output_20;
input 	temp_memtoreg_0;
input 	temp_memtoreg_1;
output 	always0;
input 	temp_regwrite1;
output 	always01;
input 	temp_branchDest_11;
input 	temp_branchDest_01;
input 	temp_branchDest_31;
input 	temp_branchDest_21;
input 	temp_branchDest_41;
output 	always02;
output 	always03;
output 	forwardb_1;
input 	temp_imemload_output_22;
input 	temp_imemload_output_21;
input 	temp_imemload_output_23;
input 	temp_imemload_output_24;
input 	temp_imemload_output_25;
output 	forwarda_1;
output 	always04;
output 	always05;
output 	always06;
output 	always07;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Equal4~0_combout ;
wire \Equal4~1_combout ;
wire \Equal1~0_combout ;
wire \always0~6_combout ;
wire \always0~5_combout ;
wire \always0~9_combout ;
wire \Equal4~2_combout ;
wire \always0~10_combout ;
wire \always0~11_combout ;
wire \Equal2~0_combout ;
wire \Equal2~1_combout ;
wire \Equal2~2_combout ;
wire \always0~4_combout ;
wire \forwarda[1]~2_combout ;
wire \always0~14_combout ;
wire \always0~15_combout ;
wire \forwarda[1]~4_combout ;
wire \Equal3~0_combout ;


// Location: LCCOMB_X59_Y41_N16
cycloneive_lcell_comb \always0~7 (
// Equation(s):
// always0 = (\Equal4~0_combout  & (\Equal4~1_combout  & (\always0~6_combout  & \always0~5_combout )))

	.dataa(\Equal4~0_combout ),
	.datab(\Equal4~1_combout ),
	.datac(\always0~6_combout ),
	.datad(\always0~5_combout ),
	.cin(gnd),
	.combout(always0),
	.cout());
// synopsys translate_off
defparam \always0~7 .lut_mask = 16'h8000;
defparam \always0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N30
cycloneive_lcell_comb \always0~8 (
// Equation(s):
// always01 = (temp_regwrite2 & ((temp_branchDest_0) # ((!temp_regwrite1) # (!\Equal1~0_combout ))))

	.dataa(temp_branchDest_0),
	.datab(\Equal1~0_combout ),
	.datac(temp_regwrite),
	.datad(temp_regwrite1),
	.cin(gnd),
	.combout(always01),
	.cout());
// synopsys translate_off
defparam \always0~8 .lut_mask = 16'hBF00;
defparam \always0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N22
cycloneive_lcell_comb \always0~12 (
// Equation(s):
// always02 = (\always0~9_combout  & (!\Equal4~2_combout  & (always01 & \always0~11_combout )))

	.dataa(\always0~9_combout ),
	.datab(\Equal4~2_combout ),
	.datac(always01),
	.datad(\always0~11_combout ),
	.cin(gnd),
	.combout(always02),
	.cout());
// synopsys translate_off
defparam \always0~12 .lut_mask = 16'h2000;
defparam \always0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N28
cycloneive_lcell_comb \always0~13 (
// Equation(s):
// always03 = (\always0~9_combout  & (!\Equal4~2_combout  & \always0~11_combout ))

	.dataa(\always0~9_combout ),
	.datab(\Equal4~2_combout ),
	.datac(gnd),
	.datad(\always0~11_combout ),
	.cin(gnd),
	.combout(always03),
	.cout());
// synopsys translate_off
defparam \always0~13 .lut_mask = 16'h2200;
defparam \always0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N22
cycloneive_lcell_comb \forwardb[1]~0 (
// Equation(s):
// forwardb_1 = (always0) # ((always01 & always03))

	.dataa(gnd),
	.datab(always0),
	.datac(always01),
	.datad(always03),
	.cin(gnd),
	.combout(forwardb_1),
	.cout());
// synopsys translate_off
defparam \forwardb[1]~0 .lut_mask = 16'hFCCC;
defparam \forwardb[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N22
cycloneive_lcell_comb \forwarda[1]~3 (
// Equation(s):
// forwarda_1 = (\Equal2~2_combout  & (((\forwarda[1]~2_combout )))) # (!\Equal2~2_combout  & (always01 & ((\forwarda[1]~4_combout ))))

	.dataa(\Equal2~2_combout ),
	.datab(always01),
	.datac(\forwarda[1]~2_combout ),
	.datad(\forwarda[1]~4_combout ),
	.cin(gnd),
	.combout(forwarda_1),
	.cout());
// synopsys translate_off
defparam \forwarda[1]~3 .lut_mask = 16'hE4A0;
defparam \forwarda[1]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N0
cycloneive_lcell_comb \always0~16 (
// Equation(s):
// always04 = (\always0~4_combout  & (!temp_memtoreg_0 & (temp_memtoreg_1 & \Equal2~2_combout )))

	.dataa(\always0~4_combout ),
	.datab(temp_memtoreg_0),
	.datac(temp_memtoreg_1),
	.datad(\Equal2~2_combout ),
	.cin(gnd),
	.combout(always04),
	.cout());
// synopsys translate_off
defparam \always0~16 .lut_mask = 16'h2000;
defparam \always0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N6
cycloneive_lcell_comb \always0~17 (
// Equation(s):
// always05 = (!\Equal2~2_combout  & (!\Equal3~0_combout  & (\always0~15_combout  & \always0~14_combout )))

	.dataa(\Equal2~2_combout ),
	.datab(\Equal3~0_combout ),
	.datac(\always0~15_combout ),
	.datad(\always0~14_combout ),
	.cin(gnd),
	.combout(always05),
	.cout());
// synopsys translate_off
defparam \always0~17 .lut_mask = 16'h1000;
defparam \always0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N24
cycloneive_lcell_comb \always0~18 (
// Equation(s):
// always06 = (\Equal4~2_combout  & (temp_regwrite1 & ((temp_branchDest_0) # (!\Equal1~0_combout ))))

	.dataa(\Equal1~0_combout ),
	.datab(\Equal4~2_combout ),
	.datac(temp_branchDest_0),
	.datad(temp_regwrite),
	.cin(gnd),
	.combout(always06),
	.cout());
// synopsys translate_off
defparam \always0~18 .lut_mask = 16'hC400;
defparam \always0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N22
cycloneive_lcell_comb \always0~19 (
// Equation(s):
// always07 = (\Equal2~2_combout  & (temp_regwrite1 & ((temp_branchDest_0) # (!\Equal1~0_combout ))))

	.dataa(\Equal2~2_combout ),
	.datab(\Equal1~0_combout ),
	.datac(temp_branchDest_0),
	.datad(temp_regwrite),
	.cin(gnd),
	.combout(always07),
	.cout());
// synopsys translate_off
defparam \always0~19 .lut_mask = 16'hA200;
defparam \always0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N30
cycloneive_lcell_comb \Equal4~0 (
// Equation(s):
// \Equal4~0_combout  = (temp_imemload_output_16 & (temp_branchDest_0 & (temp_branchDest_1 $ (!temp_imemload_output_17)))) # (!temp_imemload_output_16 & (!temp_branchDest_0 & (temp_branchDest_1 $ (!temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(temp_branchDest_1),
	.datac(temp_branchDest_0),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~0 .lut_mask = 16'h8421;
defparam \Equal4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N0
cycloneive_lcell_comb \Equal4~1 (
// Equation(s):
// \Equal4~1_combout  = (temp_branchDest_2 & (temp_imemload_output_18 & (temp_branchDest_3 $ (!temp_imemload_output_19)))) # (!temp_branchDest_2 & (!temp_imemload_output_18 & (temp_branchDest_3 $ (!temp_imemload_output_19))))

	.dataa(temp_branchDest_2),
	.datab(temp_imemload_output_18),
	.datac(temp_branchDest_3),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Equal4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~1 .lut_mask = 16'h9009;
defparam \Equal4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N2
cycloneive_lcell_comb \Equal1~0 (
// Equation(s):
// \Equal1~0_combout  = (!temp_branchDest_2 & (!temp_branchDest_3 & (!temp_branchDest_4 & !temp_branchDest_1)))

	.dataa(temp_branchDest_2),
	.datab(temp_branchDest_3),
	.datac(temp_branchDest_4),
	.datad(temp_branchDest_1),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h0001;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N26
cycloneive_lcell_comb \always0~6 (
// Equation(s):
// \always0~6_combout  = (temp_memtoreg_1 & ((temp_branchDest_0) # (!\Equal1~0_combout )))

	.dataa(gnd),
	.datab(\Equal1~0_combout ),
	.datac(temp_branchDest_0),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(\always0~6_combout ),
	.cout());
// synopsys translate_off
defparam \always0~6 .lut_mask = 16'hF300;
defparam \always0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N12
cycloneive_lcell_comb \always0~5 (
// Equation(s):
// \always0~5_combout  = (!temp_memtoreg_0 & (temp_regwrite1 & (temp_imemload_output_20 $ (!temp_branchDest_4))))

	.dataa(temp_imemload_output_20),
	.datab(temp_branchDest_4),
	.datac(temp_memtoreg_0),
	.datad(temp_regwrite),
	.cin(gnd),
	.combout(\always0~5_combout ),
	.cout());
// synopsys translate_off
defparam \always0~5 .lut_mask = 16'h0900;
defparam \always0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N24
cycloneive_lcell_comb \always0~9 (
// Equation(s):
// \always0~9_combout  = (temp_branchDest_01 & (temp_imemload_output_16 & (temp_imemload_output_17 $ (!temp_branchDest_11)))) # (!temp_branchDest_01 & (!temp_imemload_output_16 & (temp_imemload_output_17 $ (!temp_branchDest_11))))

	.dataa(temp_branchDest_01),
	.datab(temp_imemload_output_17),
	.datac(temp_branchDest_11),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\always0~9_combout ),
	.cout());
// synopsys translate_off
defparam \always0~9 .lut_mask = 16'h8241;
defparam \always0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N18
cycloneive_lcell_comb \Equal4~2 (
// Equation(s):
// \Equal4~2_combout  = (\Equal4~0_combout  & (\Equal4~1_combout  & (temp_imemload_output_20 $ (!temp_branchDest_4))))

	.dataa(temp_imemload_output_20),
	.datab(temp_branchDest_4),
	.datac(\Equal4~0_combout ),
	.datad(\Equal4~1_combout ),
	.cin(gnd),
	.combout(\Equal4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~2 .lut_mask = 16'h9000;
defparam \Equal4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N18
cycloneive_lcell_comb \always0~10 (
// Equation(s):
// \always0~10_combout  = (temp_imemload_output_18 & (temp_branchDest_21 & (temp_branchDest_31 $ (!temp_imemload_output_19)))) # (!temp_imemload_output_18 & (!temp_branchDest_21 & (temp_branchDest_31 $ (!temp_imemload_output_19))))

	.dataa(temp_imemload_output_18),
	.datab(temp_branchDest_31),
	.datac(temp_branchDest_21),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\always0~10_combout ),
	.cout());
// synopsys translate_off
defparam \always0~10 .lut_mask = 16'h8421;
defparam \always0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N6
cycloneive_lcell_comb \always0~11 (
// Equation(s):
// \always0~11_combout  = (\always0~10_combout  & (temp_branchDest_41 $ (!temp_imemload_output_20)))

	.dataa(temp_branchDest_41),
	.datab(temp_imemload_output_20),
	.datac(gnd),
	.datad(\always0~10_combout ),
	.cin(gnd),
	.combout(\always0~11_combout ),
	.cout());
// synopsys translate_off
defparam \always0~11 .lut_mask = 16'h9900;
defparam \always0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N2
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = (temp_branchDest_0 & (temp_imemload_output_21 & (temp_branchDest_1 $ (!temp_imemload_output_22)))) # (!temp_branchDest_0 & (!temp_imemload_output_21 & (temp_branchDest_1 $ (!temp_imemload_output_22))))

	.dataa(temp_branchDest_0),
	.datab(temp_imemload_output_21),
	.datac(temp_branchDest_1),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h9009;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N26
cycloneive_lcell_comb \Equal2~1 (
// Equation(s):
// \Equal2~1_combout  = (temp_branchDest_3 & (temp_imemload_output_24 & (temp_branchDest_2 $ (!temp_imemload_output_23)))) # (!temp_branchDest_3 & (!temp_imemload_output_24 & (temp_branchDest_2 $ (!temp_imemload_output_23))))

	.dataa(temp_branchDest_3),
	.datab(temp_imemload_output_24),
	.datac(temp_branchDest_2),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~1 .lut_mask = 16'h9009;
defparam \Equal2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N18
cycloneive_lcell_comb \Equal2~2 (
// Equation(s):
// \Equal2~2_combout  = (\Equal2~0_combout  & (\Equal2~1_combout  & (temp_branchDest_4 $ (!temp_imemload_output_25))))

	.dataa(temp_branchDest_4),
	.datab(\Equal2~0_combout ),
	.datac(\Equal2~1_combout ),
	.datad(temp_imemload_output_25),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~2 .lut_mask = 16'h8040;
defparam \Equal2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N20
cycloneive_lcell_comb \always0~4 (
// Equation(s):
// \always0~4_combout  = (temp_regwrite1 & ((temp_branchDest_0) # (!\Equal1~0_combout )))

	.dataa(gnd),
	.datab(\Equal1~0_combout ),
	.datac(temp_branchDest_0),
	.datad(temp_regwrite),
	.cin(gnd),
	.combout(\always0~4_combout ),
	.cout());
// synopsys translate_off
defparam \always0~4 .lut_mask = 16'hF300;
defparam \always0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N8
cycloneive_lcell_comb \forwarda[1]~2 (
// Equation(s):
// \forwarda[1]~2_combout  = (temp_memtoreg_1 & (\always0~4_combout  & !temp_memtoreg_0))

	.dataa(temp_memtoreg_1),
	.datab(gnd),
	.datac(\always0~4_combout ),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(\forwarda[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \forwarda[1]~2 .lut_mask = 16'h00A0;
defparam \forwarda[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N10
cycloneive_lcell_comb \always0~14 (
// Equation(s):
// \always0~14_combout  = (temp_imemload_output_22 & (temp_branchDest_11 & (temp_branchDest_01 $ (!temp_imemload_output_21)))) # (!temp_imemload_output_22 & (!temp_branchDest_11 & (temp_branchDest_01 $ (!temp_imemload_output_21))))

	.dataa(temp_imemload_output_22),
	.datab(temp_branchDest_11),
	.datac(temp_branchDest_01),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\always0~14_combout ),
	.cout());
// synopsys translate_off
defparam \always0~14 .lut_mask = 16'h9009;
defparam \always0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N8
cycloneive_lcell_comb \always0~15 (
// Equation(s):
// \always0~15_combout  = (temp_branchDest_31 & (temp_imemload_output_24 & (temp_branchDest_21 $ (!temp_imemload_output_23)))) # (!temp_branchDest_31 & (!temp_imemload_output_24 & (temp_branchDest_21 $ (!temp_imemload_output_23))))

	.dataa(temp_branchDest_31),
	.datab(temp_imemload_output_24),
	.datac(temp_branchDest_21),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\always0~15_combout ),
	.cout());
// synopsys translate_off
defparam \always0~15 .lut_mask = 16'h9009;
defparam \always0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N10
cycloneive_lcell_comb \forwarda[1]~4 (
// Equation(s):
// \forwarda[1]~4_combout  = (\always0~14_combout  & (\always0~15_combout  & (temp_imemload_output_25 $ (!temp_branchDest_41))))

	.dataa(\always0~14_combout ),
	.datab(temp_imemload_output_25),
	.datac(\always0~15_combout ),
	.datad(temp_branchDest_41),
	.cin(gnd),
	.combout(\forwarda[1]~4_combout ),
	.cout());
// synopsys translate_off
defparam \forwarda[1]~4 .lut_mask = 16'h8020;
defparam \forwarda[1]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N20
cycloneive_lcell_comb \Equal3~0 (
// Equation(s):
// \Equal3~0_combout  = temp_branchDest_41 $ (temp_imemload_output_25)

	.dataa(gnd),
	.datab(temp_branchDest_41),
	.datac(gnd),
	.datad(temp_imemload_output_25),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~0 .lut_mask = 16'h33CC;
defparam \Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module hazard_unit (
	temp_zeroFlag,
	temp_dmemWEN,
	temp_dmemREN,
	always1,
	temp_halt_out,
	temp_imemload_output_17,
	temp_imemload_output_16,
	temp_imemload_output_18,
	temp_imemload_output_19,
	temp_imemload_output_20,
	temp_iMemLoad_0,
	temp_iMemLoad_1,
	temp_iMemLoad_4,
	temp_iMemLoad_3,
	temp_iMemLoad_2,
	temp_iMemLoad_5,
	temp_iMemLoad_31,
	temp_iMemLoad_30,
	temp_iMemLoad_29,
	ex_mem_flush,
	temp_iMemLoad_27,
	temp_iMemLoad_26,
	temp_iMemLoad_28,
	ex_mem_flush1,
	temp_branchSelect,
	ex_mem_flush2,
	ex_mem_flush3,
	id_ex_wen,
	ccifiwait_0,
	temp_request_dmemREN_output,
	temp_imemload_output_171,
	temp_imemload_output_161,
	temp_imemload_output_191,
	temp_imemload_output_181,
	temp_imemload_output_201,
	temp_imemload_output_22,
	temp_imemload_output_21,
	temp_imemload_output_24,
	temp_imemload_output_23,
	temp_imemload_output_25,
	use_after_load,
	pc_wen,
	id_ex_flush1,
	pc_wen1,
	devpor,
	devclrn,
	devoe);
input 	temp_zeroFlag;
input 	temp_dmemWEN;
input 	temp_dmemREN;
input 	always1;
input 	temp_halt_out;
input 	temp_imemload_output_17;
input 	temp_imemload_output_16;
input 	temp_imemload_output_18;
input 	temp_imemload_output_19;
input 	temp_imemload_output_20;
input 	temp_iMemLoad_0;
input 	temp_iMemLoad_1;
input 	temp_iMemLoad_4;
input 	temp_iMemLoad_3;
input 	temp_iMemLoad_2;
input 	temp_iMemLoad_5;
input 	temp_iMemLoad_31;
input 	temp_iMemLoad_30;
input 	temp_iMemLoad_29;
output 	ex_mem_flush;
input 	temp_iMemLoad_27;
input 	temp_iMemLoad_26;
input 	temp_iMemLoad_28;
output 	ex_mem_flush1;
input 	temp_branchSelect;
output 	ex_mem_flush2;
output 	ex_mem_flush3;
output 	id_ex_wen;
input 	ccifiwait_0;
input 	temp_request_dmemREN_output;
input 	temp_imemload_output_171;
input 	temp_imemload_output_161;
input 	temp_imemload_output_191;
input 	temp_imemload_output_181;
input 	temp_imemload_output_201;
input 	temp_imemload_output_22;
input 	temp_imemload_output_21;
input 	temp_imemload_output_24;
input 	temp_imemload_output_23;
input 	temp_imemload_output_25;
output 	use_after_load;
output 	pc_wen;
output 	id_ex_flush1;
output 	pc_wen1;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \ex_mem_flush~1_combout ;
wire \ex_mem_flush~2_combout ;
wire \use_after_load~1_combout ;
wire \use_after_load~0_combout ;
wire \use_after_load~2_combout ;
wire \use_after_load~4_combout ;
wire \use_after_load~3_combout ;
wire \use_after_load~5_combout ;
wire \pc_wen~4_combout ;


// Location: LCCOMB_X62_Y38_N18
cycloneive_lcell_comb \ex_mem_flush~0 (
// Equation(s):
// ex_mem_flush = (!temp_iMemLoad_31 & (!temp_iMemLoad_30 & !temp_iMemLoad_29))

	.dataa(temp_iMemLoad_31),
	.datab(temp_iMemLoad_30),
	.datac(gnd),
	.datad(temp_iMemLoad_29),
	.cin(gnd),
	.combout(ex_mem_flush),
	.cout());
// synopsys translate_off
defparam \ex_mem_flush~0 .lut_mask = 16'h0011;
defparam \ex_mem_flush~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N22
cycloneive_lcell_comb \ex_mem_flush~3 (
// Equation(s):
// ex_mem_flush1 = (!temp_iMemLoad_28 & ((temp_iMemLoad_27) # ((\ex_mem_flush~1_combout  & \ex_mem_flush~2_combout ))))

	.dataa(\ex_mem_flush~1_combout ),
	.datab(temp_iMemLoad_28),
	.datac(\ex_mem_flush~2_combout ),
	.datad(temp_iMemLoad_27),
	.cin(gnd),
	.combout(ex_mem_flush1),
	.cout());
// synopsys translate_off
defparam \ex_mem_flush~3 .lut_mask = 16'h3320;
defparam \ex_mem_flush~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N20
cycloneive_lcell_comb \ex_mem_flush~4 (
// Equation(s):
// ex_mem_flush2 = (temp_iMemLoad_28 & (!temp_iMemLoad_27 & (temp_zeroFlag1 $ (!temp_branchSelect1))))

	.dataa(temp_zeroFlag),
	.datab(temp_iMemLoad_28),
	.datac(temp_branchSelect),
	.datad(temp_iMemLoad_27),
	.cin(gnd),
	.combout(ex_mem_flush2),
	.cout());
// synopsys translate_off
defparam \ex_mem_flush~4 .lut_mask = 16'h0084;
defparam \ex_mem_flush~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N4
cycloneive_lcell_comb \ex_mem_flush~5 (
// Equation(s):
// ex_mem_flush3 = (ex_mem_flush & ((ex_mem_flush2) # (ex_mem_flush1)))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ex_mem_flush2),
	.datad(ex_mem_flush1),
	.cin(gnd),
	.combout(ex_mem_flush3),
	.cout());
// synopsys translate_off
defparam \ex_mem_flush~5 .lut_mask = 16'hCCC0;
defparam \ex_mem_flush~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N26
cycloneive_lcell_comb \id_ex_wen~0 (
// Equation(s):
// id_ex_wen = (!temp_halt_out1 & ((always1) # ((!temp_dmemREN1 & !temp_dmemWEN1))))

	.dataa(temp_dmemREN),
	.datab(temp_dmemWEN),
	.datac(always1),
	.datad(temp_halt_out),
	.cin(gnd),
	.combout(id_ex_wen),
	.cout());
// synopsys translate_off
defparam \id_ex_wen~0 .lut_mask = 16'h00F1;
defparam \id_ex_wen~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N24
cycloneive_lcell_comb \use_after_load~6 (
// Equation(s):
// use_after_load = (temp_request_dmemREN_output1 & ((\use_after_load~2_combout ) # (\use_after_load~5_combout )))

	.dataa(gnd),
	.datab(\use_after_load~2_combout ),
	.datac(\use_after_load~5_combout ),
	.datad(temp_request_dmemREN_output),
	.cin(gnd),
	.combout(use_after_load),
	.cout());
// synopsys translate_off
defparam \use_after_load~6 .lut_mask = 16'hFC00;
defparam \use_after_load~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N6
cycloneive_lcell_comb \pc_wen~2 (
// Equation(s):
// pc_wen = (id_ex_wen & (!use_after_load & ((ex_mem_flush3) # (!ccifiwait_0))))

	.dataa(id_ex_wen),
	.datab(use_after_load),
	.datac(ccifiwait_0),
	.datad(ex_mem_flush3),
	.cin(gnd),
	.combout(pc_wen),
	.cout());
// synopsys translate_off
defparam \pc_wen~2 .lut_mask = 16'h2202;
defparam \pc_wen~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N14
cycloneive_lcell_comb id_ex_flush(
// Equation(s):
// id_ex_flush1 = (ex_mem_flush3) # ((temp_request_dmemREN_output1 & ((\use_after_load~5_combout ) # (\use_after_load~2_combout ))))

	.dataa(\use_after_load~5_combout ),
	.datab(\use_after_load~2_combout ),
	.datac(ex_mem_flush3),
	.datad(temp_request_dmemREN_output),
	.cin(gnd),
	.combout(id_ex_flush1),
	.cout());
// synopsys translate_off
defparam id_ex_flush.lut_mask = 16'hFEF0;
defparam id_ex_flush.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N20
cycloneive_lcell_comb \pc_wen~3 (
// Equation(s):
// pc_wen1 = (\pc_wen~4_combout  & ((always1) # ((!temp_dmemREN1 & !temp_dmemWEN1))))

	.dataa(temp_dmemREN),
	.datab(temp_dmemWEN),
	.datac(always1),
	.datad(\pc_wen~4_combout ),
	.cin(gnd),
	.combout(pc_wen1),
	.cout());
// synopsys translate_off
defparam \pc_wen~3 .lut_mask = 16'hF100;
defparam \pc_wen~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N12
cycloneive_lcell_comb \ex_mem_flush~1 (
// Equation(s):
// \ex_mem_flush~1_combout  = (!temp_iMemLoad_4 & (!temp_iMemLoad_26 & (!temp_iMemLoad_5 & temp_iMemLoad_3)))

	.dataa(temp_iMemLoad_4),
	.datab(temp_iMemLoad_26),
	.datac(temp_iMemLoad_5),
	.datad(temp_iMemLoad_3),
	.cin(gnd),
	.combout(\ex_mem_flush~1_combout ),
	.cout());
// synopsys translate_off
defparam \ex_mem_flush~1 .lut_mask = 16'h0100;
defparam \ex_mem_flush~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N14
cycloneive_lcell_comb \ex_mem_flush~2 (
// Equation(s):
// \ex_mem_flush~2_combout  = (!temp_iMemLoad_0 & (!temp_iMemLoad_2 & !temp_iMemLoad_1))

	.dataa(temp_iMemLoad_0),
	.datab(temp_iMemLoad_2),
	.datac(gnd),
	.datad(temp_iMemLoad_1),
	.cin(gnd),
	.combout(\ex_mem_flush~2_combout ),
	.cout());
// synopsys translate_off
defparam \ex_mem_flush~2 .lut_mask = 16'h0011;
defparam \ex_mem_flush~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N2
cycloneive_lcell_comb \use_after_load~1 (
// Equation(s):
// \use_after_load~1_combout  = (temp_imemload_output_19 & (temp_imemload_output_19 & (temp_imemload_output_18 $ (!temp_imemload_output_18)))) # (!temp_imemload_output_19 & (!temp_imemload_output_19 & (temp_imemload_output_18 $ (!temp_imemload_output_18))))

	.dataa(temp_imemload_output_191),
	.datab(temp_imemload_output_18),
	.datac(temp_imemload_output_181),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\use_after_load~1_combout ),
	.cout());
// synopsys translate_off
defparam \use_after_load~1 .lut_mask = 16'h8241;
defparam \use_after_load~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N6
cycloneive_lcell_comb \use_after_load~0 (
// Equation(s):
// \use_after_load~0_combout  = (temp_imemload_output_16 & (temp_imemload_output_16 & (temp_imemload_output_17 $ (!temp_imemload_output_17)))) # (!temp_imemload_output_16 & (!temp_imemload_output_16 & (temp_imemload_output_17 $ (!temp_imemload_output_17))))

	.dataa(temp_imemload_output_161),
	.datab(temp_imemload_output_17),
	.datac(temp_imemload_output_171),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\use_after_load~0_combout ),
	.cout());
// synopsys translate_off
defparam \use_after_load~0 .lut_mask = 16'h8241;
defparam \use_after_load~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N8
cycloneive_lcell_comb \use_after_load~2 (
// Equation(s):
// \use_after_load~2_combout  = (\use_after_load~1_combout  & (\use_after_load~0_combout  & (temp_imemload_output_20 $ (!temp_imemload_output_20))))

	.dataa(temp_imemload_output_20),
	.datab(temp_imemload_output_201),
	.datac(\use_after_load~1_combout ),
	.datad(\use_after_load~0_combout ),
	.cin(gnd),
	.combout(\use_after_load~2_combout ),
	.cout());
// synopsys translate_off
defparam \use_after_load~2 .lut_mask = 16'h9000;
defparam \use_after_load~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N26
cycloneive_lcell_comb \use_after_load~4 (
// Equation(s):
// \use_after_load~4_combout  = (temp_imemload_output_18 & (temp_imemload_output_23 & (temp_imemload_output_24 $ (!temp_imemload_output_19)))) # (!temp_imemload_output_18 & (!temp_imemload_output_23 & (temp_imemload_output_24 $ (!temp_imemload_output_19))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_24),
	.datac(temp_imemload_output_19),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\use_after_load~4_combout ),
	.cout());
// synopsys translate_off
defparam \use_after_load~4 .lut_mask = 16'h8241;
defparam \use_after_load~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N4
cycloneive_lcell_comb \use_after_load~3 (
// Equation(s):
// \use_after_load~3_combout  = (temp_imemload_output_21 & (temp_imemload_output_16 & (temp_imemload_output_17 $ (!temp_imemload_output_22)))) # (!temp_imemload_output_21 & (!temp_imemload_output_16 & (temp_imemload_output_17 $ (!temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_17),
	.datac(temp_imemload_output_22),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\use_after_load~3_combout ),
	.cout());
// synopsys translate_off
defparam \use_after_load~3 .lut_mask = 16'h8241;
defparam \use_after_load~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N22
cycloneive_lcell_comb \use_after_load~5 (
// Equation(s):
// \use_after_load~5_combout  = (\use_after_load~4_combout  & (\use_after_load~3_combout  & (temp_imemload_output_20 $ (!temp_imemload_output_25))))

	.dataa(temp_imemload_output_20),
	.datab(\use_after_load~4_combout ),
	.datac(temp_imemload_output_25),
	.datad(\use_after_load~3_combout ),
	.cin(gnd),
	.combout(\use_after_load~5_combout ),
	.cout());
// synopsys translate_off
defparam \use_after_load~5 .lut_mask = 16'h8400;
defparam \use_after_load~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N4
cycloneive_lcell_comb \pc_wen~4 (
// Equation(s):
// \pc_wen~4_combout  = (!temp_halt_out1 & (((!\use_after_load~2_combout  & !\use_after_load~5_combout )) # (!temp_request_dmemREN_output1)))

	.dataa(temp_halt_out),
	.datab(\use_after_load~2_combout ),
	.datac(\use_after_load~5_combout ),
	.datad(temp_request_dmemREN_output),
	.cin(gnd),
	.combout(\pc_wen~4_combout ),
	.cout());
// synopsys translate_off
defparam \pc_wen~4 .lut_mask = 16'h0155;
defparam \pc_wen~4 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module id_ex_latch (
	temp_signzerovalue_output_16,
	temp_halt_out_output1,
	temp_ALUop_output_0,
	temp_imemload_output_1,
	temp_imemload_output_7,
	temp_ALUsrc_output_1,
	temp_ALUsrc_output_0,
	temp_rdat_two_output_1,
	temp_imemload_output_17,
	temp_imemload_output_16,
	temp_imemload_output_18,
	temp_imemload_output_19,
	temp_imemload_output_20,
	temp_imemload_output_22,
	temp_imemload_output_21,
	temp_imemload_output_23,
	temp_imemload_output_24,
	temp_imemload_output_25,
	temp_rdat_one_output_1,
	temp_ALUop_output_1,
	temp_imemload_output_0,
	temp_imemload_output_6,
	temp_rdat_two_output_0,
	temp_rdat_one_output_0,
	temp_rdat_one_output_2,
	temp_rdat_one_output_4,
	temp_rdat_one_output_3,
	temp_imemload_output_2,
	temp_imemload_output_8,
	temp_rdat_two_output_2,
	temp_rdat_one_output_8,
	temp_rdat_one_output_7,
	temp_rdat_one_output_6,
	temp_rdat_one_output_5,
	temp_imemload_output_3,
	temp_imemload_output_9,
	temp_rdat_two_output_3,
	temp_rdat_one_output_16,
	temp_rdat_one_output_14,
	temp_rdat_one_output_15,
	temp_rdat_one_output_13,
	temp_rdat_one_output_12,
	temp_rdat_one_output_10,
	temp_rdat_one_output_11,
	temp_rdat_one_output_9,
	temp_imemload_output_4,
	temp_imemload_output_10,
	temp_rdat_two_output_4,
	temp_rdat_one_output_31,
	temp_rdat_one_output_30,
	temp_rdat_one_output_29,
	temp_rdat_one_output_26,
	temp_rdat_one_output_25,
	temp_rdat_one_output_28,
	temp_rdat_one_output_27,
	temp_rdat_one_output_17,
	temp_rdat_one_output_20,
	temp_rdat_one_output_19,
	temp_rdat_one_output_18,
	temp_rdat_one_output_24,
	temp_rdat_one_output_23,
	temp_rdat_one_output_22,
	temp_rdat_one_output_21,
	temp_rdat_two_output_15,
	temp_imemload_output_15,
	temp_rdat_two_output_12,
	temp_imemload_output_12,
	temp_rdat_two_output_27,
	temp_rdat_two_output_18,
	temp_rdat_two_output_17,
	temp_rdat_two_output_16,
	temp_rdat_two_output_31,
	temp_rdat_two_output_30,
	temp_rdat_two_output_29,
	temp_rdat_two_output_28,
	temp_rdat_two_output_26,
	temp_rdat_two_output_25,
	temp_rdat_two_output_24,
	temp_rdat_two_output_23,
	temp_rdat_two_output_22,
	temp_rdat_two_output_21,
	temp_rdat_two_output_20,
	temp_rdat_two_output_19,
	temp_imemload_output_14,
	temp_rdat_two_output_10,
	temp_rdat_two_output_14,
	temp_rdat_two_output_9,
	temp_rdat_two_output_8,
	temp_rdat_two_output_7,
	temp_rdat_two_output_6,
	temp_rdat_two_output_5,
	temp_imemload_output_5,
	temp_rdat_two_output_13,
	temp_imemload_output_13,
	temp_rdat_two_output_11,
	temp_imemload_output_11,
	temp_ALUop_output_2,
	temp_ALUop_output_3,
	ex_mem_flush,
	wen,
	temp_request_dmemREN_output1,
	temp_imemload_output_171,
	temp_imemload_output_161,
	temp_imemload_output_191,
	temp_imemload_output_181,
	temp_imemload_output_201,
	temp_imemload_output_221,
	temp_imemload_output_211,
	temp_imemload_output_241,
	temp_imemload_output_231,
	temp_imemload_output_251,
	use_after_load,
	temp_request_dmemWEN_output1,
	temp_imemload_output_29,
	temp_imemload_output_31,
	temp_imemload_output_30,
	temp_imemload_output_28,
	Equal3,
	temp_imemload_output_27,
	temp_imemload_output_26,
	temp_branch_output1,
	temp_imemload_output_01,
	temp_imemload_output_210,
	temp_imemload_output_32,
	temp_imemload_output_51,
	Equal31,
	temp_imemload_output_151,
	temp_imemload_output_141,
	temp_imemload_output_131,
	temp_imemload_output_121,
	temp_imemload_output_111,
	temp_imemload_output_101,
	temp_imemload_output_91,
	temp_imemload_output_81,
	temp_imemload_output_71,
	temp_imemload_output_61,
	temp_imemload_output_110,
	temp_imemload_output_41,
	Equal32,
	extended_imm_16,
	WideOr8,
	WideOr2,
	id_ex_flush,
	WideOr4,
	temp_ALUsrc_output,
	Mux62,
	Mux621,
	temp_regwrite_output1,
	temp_regdst_output_1,
	temp_regdst_output_0,
	temp_memtoreg_output_0,
	temp_memtoreg_output_1,
	Mux30,
	Mux301,
	WideOr7,
	WideOr1,
	Mux63,
	Mux631,
	Mux31,
	Mux311,
	Mux29,
	Mux291,
	Mux27,
	Mux271,
	Mux28,
	Mux281,
	Mux61,
	Mux611,
	Mux23,
	Mux231,
	Mux24,
	Mux241,
	Mux25,
	Mux251,
	Mux26,
	Mux261,
	Mux60,
	Mux601,
	Mux15,
	Mux151,
	Mux17,
	Mux171,
	Mux16,
	Mux161,
	Mux18,
	Mux181,
	Mux19,
	Mux191,
	Mux21,
	Mux211,
	Mux20,
	Mux201,
	Mux22,
	Mux221,
	Mux59,
	Mux591,
	Mux0,
	Mux01,
	Mux1,
	Mux11,
	Mux2,
	Mux210,
	Mux5,
	Mux51,
	Mux6,
	Mux64,
	Mux3,
	Mux32,
	Mux4,
	Mux41,
	Mux14,
	Mux141,
	Mux111,
	Mux112,
	Mux12,
	Mux121,
	Mux13,
	Mux131,
	Mux7,
	Mux71,
	Mux8,
	Mux81,
	Mux9,
	Mux91,
	Mux10,
	Mux101,
	Mux48,
	Mux481,
	Mux511,
	Mux512,
	Mux36,
	Mux361,
	extended_imm_161,
	Mux45,
	Mux451,
	Mux46,
	Mux461,
	Mux47,
	Mux471,
	Mux321,
	Mux322,
	Mux33,
	Mux331,
	Mux34,
	Mux341,
	Mux35,
	Mux351,
	Mux37,
	Mux371,
	Mux38,
	Mux381,
	Mux39,
	Mux391,
	Mux40,
	Mux401,
	Mux411,
	Mux412,
	Mux42,
	Mux421,
	Mux43,
	Mux431,
	Mux44,
	Mux441,
	Mux53,
	Mux531,
	Mux49,
	Mux491,
	Mux54,
	Mux541,
	Mux55,
	Mux551,
	Mux56,
	Mux561,
	Mux57,
	Mux571,
	Mux58,
	Mux581,
	Mux50,
	Mux501,
	Mux52,
	Mux521,
	WideOr6,
	WideOr0,
	halt_out,
	temp_imemload_output_311,
	temp_imemload_output_301,
	temp_imemload_output_291,
	temp_imemload_output_271,
	temp_imemload_output_261,
	temp_imemload_output_281,
	temp_branch_output2,
	temp_NPC_output_1,
	temp_pcselect_output_1,
	temp_pcselect_output_0,
	temp_NPC_output_0,
	temp_NPC_output_2,
	temp_NPC_output_3,
	temp_NPC_output_5,
	temp_NPC_output_4,
	temp_NPC_output_7,
	temp_NPC_output_6,
	temp_NPC_output_9,
	temp_NPC_output_8,
	temp_NPC_output_11,
	temp_NPC_output_10,
	temp_NPC_output_13,
	temp_NPC_output_12,
	temp_NPC_output_15,
	temp_NPC_output_14,
	temp_NPC_output_17,
	temp_NPC_output_16,
	temp_NPC_output_19,
	temp_NPC_output_18,
	temp_NPC_output_20,
	temp_NPC_output_21,
	temp_NPC_output_23,
	temp_NPC_output_22,
	temp_NPC_output_25,
	temp_NPC_output_24,
	temp_NPC_output_26,
	temp_NPC_output_27,
	temp_NPC_output_29,
	temp_NPC_output_28,
	temp_NPC_output_31,
	temp_NPC_output_30,
	halt_out1,
	WideOr3,
	WideOr10,
	memtoreg,
	temp_NPC_output_110,
	WideOr9,
	temp_NPC_output_01,
	temp_NPC_output_210,
	temp_NPC_output_32,
	temp_NPC_output_51,
	temp_NPC_output_41,
	temp_NPC_output_71,
	temp_NPC_output_61,
	temp_NPC_output_91,
	temp_NPC_output_81,
	temp_NPC_output_111,
	temp_NPC_output_101,
	temp_NPC_output_131,
	temp_NPC_output_121,
	temp_NPC_output_151,
	temp_NPC_output_141,
	temp_NPC_output_171,
	temp_NPC_output_161,
	temp_NPC_output_191,
	temp_NPC_output_181,
	temp_NPC_output_201,
	temp_NPC_output_211,
	temp_NPC_output_231,
	temp_NPC_output_221,
	temp_NPC_output_251,
	temp_NPC_output_241,
	temp_NPC_output_261,
	temp_NPC_output_271,
	temp_NPC_output_291,
	temp_NPC_output_281,
	temp_NPC_output_311,
	temp_NPC_output_301,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	temp_signzerovalue_output_16;
output 	temp_halt_out_output1;
output 	temp_ALUop_output_0;
output 	temp_imemload_output_1;
output 	temp_imemload_output_7;
output 	temp_ALUsrc_output_1;
output 	temp_ALUsrc_output_0;
output 	temp_rdat_two_output_1;
output 	temp_imemload_output_17;
output 	temp_imemload_output_16;
output 	temp_imemload_output_18;
output 	temp_imemload_output_19;
output 	temp_imemload_output_20;
output 	temp_imemload_output_22;
output 	temp_imemload_output_21;
output 	temp_imemload_output_23;
output 	temp_imemload_output_24;
output 	temp_imemload_output_25;
output 	temp_rdat_one_output_1;
output 	temp_ALUop_output_1;
output 	temp_imemload_output_0;
output 	temp_imemload_output_6;
output 	temp_rdat_two_output_0;
output 	temp_rdat_one_output_0;
output 	temp_rdat_one_output_2;
output 	temp_rdat_one_output_4;
output 	temp_rdat_one_output_3;
output 	temp_imemload_output_2;
output 	temp_imemload_output_8;
output 	temp_rdat_two_output_2;
output 	temp_rdat_one_output_8;
output 	temp_rdat_one_output_7;
output 	temp_rdat_one_output_6;
output 	temp_rdat_one_output_5;
output 	temp_imemload_output_3;
output 	temp_imemload_output_9;
output 	temp_rdat_two_output_3;
output 	temp_rdat_one_output_16;
output 	temp_rdat_one_output_14;
output 	temp_rdat_one_output_15;
output 	temp_rdat_one_output_13;
output 	temp_rdat_one_output_12;
output 	temp_rdat_one_output_10;
output 	temp_rdat_one_output_11;
output 	temp_rdat_one_output_9;
output 	temp_imemload_output_4;
output 	temp_imemload_output_10;
output 	temp_rdat_two_output_4;
output 	temp_rdat_one_output_31;
output 	temp_rdat_one_output_30;
output 	temp_rdat_one_output_29;
output 	temp_rdat_one_output_26;
output 	temp_rdat_one_output_25;
output 	temp_rdat_one_output_28;
output 	temp_rdat_one_output_27;
output 	temp_rdat_one_output_17;
output 	temp_rdat_one_output_20;
output 	temp_rdat_one_output_19;
output 	temp_rdat_one_output_18;
output 	temp_rdat_one_output_24;
output 	temp_rdat_one_output_23;
output 	temp_rdat_one_output_22;
output 	temp_rdat_one_output_21;
output 	temp_rdat_two_output_15;
output 	temp_imemload_output_15;
output 	temp_rdat_two_output_12;
output 	temp_imemload_output_12;
output 	temp_rdat_two_output_27;
output 	temp_rdat_two_output_18;
output 	temp_rdat_two_output_17;
output 	temp_rdat_two_output_16;
output 	temp_rdat_two_output_31;
output 	temp_rdat_two_output_30;
output 	temp_rdat_two_output_29;
output 	temp_rdat_two_output_28;
output 	temp_rdat_two_output_26;
output 	temp_rdat_two_output_25;
output 	temp_rdat_two_output_24;
output 	temp_rdat_two_output_23;
output 	temp_rdat_two_output_22;
output 	temp_rdat_two_output_21;
output 	temp_rdat_two_output_20;
output 	temp_rdat_two_output_19;
output 	temp_imemload_output_14;
output 	temp_rdat_two_output_10;
output 	temp_rdat_two_output_14;
output 	temp_rdat_two_output_9;
output 	temp_rdat_two_output_8;
output 	temp_rdat_two_output_7;
output 	temp_rdat_two_output_6;
output 	temp_rdat_two_output_5;
output 	temp_imemload_output_5;
output 	temp_rdat_two_output_13;
output 	temp_imemload_output_13;
output 	temp_rdat_two_output_11;
output 	temp_imemload_output_11;
output 	temp_ALUop_output_2;
output 	temp_ALUop_output_3;
input 	ex_mem_flush;
input 	wen;
output 	temp_request_dmemREN_output1;
input 	temp_imemload_output_171;
input 	temp_imemload_output_161;
input 	temp_imemload_output_191;
input 	temp_imemload_output_181;
input 	temp_imemload_output_201;
input 	temp_imemload_output_221;
input 	temp_imemload_output_211;
input 	temp_imemload_output_241;
input 	temp_imemload_output_231;
input 	temp_imemload_output_251;
input 	use_after_load;
output 	temp_request_dmemWEN_output1;
input 	temp_imemload_output_29;
input 	temp_imemload_output_31;
input 	temp_imemload_output_30;
input 	temp_imemload_output_28;
input 	Equal3;
input 	temp_imemload_output_27;
input 	temp_imemload_output_26;
output 	temp_branch_output1;
input 	temp_imemload_output_01;
input 	temp_imemload_output_210;
input 	temp_imemload_output_32;
input 	temp_imemload_output_51;
input 	Equal31;
input 	temp_imemload_output_151;
input 	temp_imemload_output_141;
input 	temp_imemload_output_131;
input 	temp_imemload_output_121;
input 	temp_imemload_output_111;
input 	temp_imemload_output_101;
input 	temp_imemload_output_91;
input 	temp_imemload_output_81;
input 	temp_imemload_output_71;
input 	temp_imemload_output_61;
input 	temp_imemload_output_110;
input 	temp_imemload_output_41;
input 	Equal32;
input 	extended_imm_16;
input 	WideOr8;
input 	WideOr2;
input 	id_ex_flush;
input 	WideOr4;
output 	temp_ALUsrc_output;
input 	Mux62;
input 	Mux621;
output 	temp_regwrite_output1;
output 	temp_regdst_output_1;
output 	temp_regdst_output_0;
output 	temp_memtoreg_output_0;
output 	temp_memtoreg_output_1;
input 	Mux30;
input 	Mux301;
input 	WideOr7;
input 	WideOr1;
input 	Mux63;
input 	Mux631;
input 	Mux31;
input 	Mux311;
input 	Mux29;
input 	Mux291;
input 	Mux27;
input 	Mux271;
input 	Mux28;
input 	Mux281;
input 	Mux61;
input 	Mux611;
input 	Mux23;
input 	Mux231;
input 	Mux24;
input 	Mux241;
input 	Mux25;
input 	Mux251;
input 	Mux26;
input 	Mux261;
input 	Mux60;
input 	Mux601;
input 	Mux15;
input 	Mux151;
input 	Mux17;
input 	Mux171;
input 	Mux16;
input 	Mux161;
input 	Mux18;
input 	Mux181;
input 	Mux19;
input 	Mux191;
input 	Mux21;
input 	Mux211;
input 	Mux20;
input 	Mux201;
input 	Mux22;
input 	Mux221;
input 	Mux59;
input 	Mux591;
input 	Mux0;
input 	Mux01;
input 	Mux1;
input 	Mux11;
input 	Mux2;
input 	Mux210;
input 	Mux5;
input 	Mux51;
input 	Mux6;
input 	Mux64;
input 	Mux3;
input 	Mux32;
input 	Mux4;
input 	Mux41;
input 	Mux14;
input 	Mux141;
input 	Mux111;
input 	Mux112;
input 	Mux12;
input 	Mux121;
input 	Mux13;
input 	Mux131;
input 	Mux7;
input 	Mux71;
input 	Mux8;
input 	Mux81;
input 	Mux9;
input 	Mux91;
input 	Mux10;
input 	Mux101;
input 	Mux48;
input 	Mux481;
input 	Mux511;
input 	Mux512;
input 	Mux36;
input 	Mux361;
input 	extended_imm_161;
input 	Mux45;
input 	Mux451;
input 	Mux46;
input 	Mux461;
input 	Mux47;
input 	Mux471;
input 	Mux321;
input 	Mux322;
input 	Mux33;
input 	Mux331;
input 	Mux34;
input 	Mux341;
input 	Mux35;
input 	Mux351;
input 	Mux37;
input 	Mux371;
input 	Mux38;
input 	Mux381;
input 	Mux39;
input 	Mux391;
input 	Mux40;
input 	Mux401;
input 	Mux411;
input 	Mux412;
input 	Mux42;
input 	Mux421;
input 	Mux43;
input 	Mux431;
input 	Mux44;
input 	Mux441;
input 	Mux53;
input 	Mux531;
input 	Mux49;
input 	Mux491;
input 	Mux54;
input 	Mux541;
input 	Mux55;
input 	Mux551;
input 	Mux56;
input 	Mux561;
input 	Mux57;
input 	Mux571;
input 	Mux58;
input 	Mux581;
input 	Mux50;
input 	Mux501;
input 	Mux52;
input 	Mux521;
input 	WideOr6;
input 	WideOr0;
input 	halt_out;
output 	temp_imemload_output_311;
output 	temp_imemload_output_301;
output 	temp_imemload_output_291;
output 	temp_imemload_output_271;
output 	temp_imemload_output_261;
output 	temp_imemload_output_281;
output 	temp_branch_output2;
output 	temp_NPC_output_1;
output 	temp_pcselect_output_1;
output 	temp_pcselect_output_0;
output 	temp_NPC_output_0;
output 	temp_NPC_output_2;
output 	temp_NPC_output_3;
output 	temp_NPC_output_5;
output 	temp_NPC_output_4;
output 	temp_NPC_output_7;
output 	temp_NPC_output_6;
output 	temp_NPC_output_9;
output 	temp_NPC_output_8;
output 	temp_NPC_output_11;
output 	temp_NPC_output_10;
output 	temp_NPC_output_13;
output 	temp_NPC_output_12;
output 	temp_NPC_output_15;
output 	temp_NPC_output_14;
output 	temp_NPC_output_17;
output 	temp_NPC_output_16;
output 	temp_NPC_output_19;
output 	temp_NPC_output_18;
output 	temp_NPC_output_20;
output 	temp_NPC_output_21;
output 	temp_NPC_output_23;
output 	temp_NPC_output_22;
output 	temp_NPC_output_25;
output 	temp_NPC_output_24;
output 	temp_NPC_output_26;
output 	temp_NPC_output_27;
output 	temp_NPC_output_29;
output 	temp_NPC_output_28;
output 	temp_NPC_output_31;
output 	temp_NPC_output_30;
input 	halt_out1;
input 	WideOr3;
input 	WideOr10;
input 	memtoreg;
input 	temp_NPC_output_110;
input 	WideOr9;
input 	temp_NPC_output_01;
input 	temp_NPC_output_210;
input 	temp_NPC_output_32;
input 	temp_NPC_output_51;
input 	temp_NPC_output_41;
input 	temp_NPC_output_71;
input 	temp_NPC_output_61;
input 	temp_NPC_output_91;
input 	temp_NPC_output_81;
input 	temp_NPC_output_111;
input 	temp_NPC_output_101;
input 	temp_NPC_output_131;
input 	temp_NPC_output_121;
input 	temp_NPC_output_151;
input 	temp_NPC_output_141;
input 	temp_NPC_output_171;
input 	temp_NPC_output_161;
input 	temp_NPC_output_191;
input 	temp_NPC_output_181;
input 	temp_NPC_output_201;
input 	temp_NPC_output_211;
input 	temp_NPC_output_231;
input 	temp_NPC_output_221;
input 	temp_NPC_output_251;
input 	temp_NPC_output_241;
input 	temp_NPC_output_261;
input 	temp_NPC_output_271;
input 	temp_NPC_output_291;
input 	temp_NPC_output_281;
input 	temp_NPC_output_311;
input 	temp_NPC_output_301;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \temp_ALUop_output~2_combout ;
wire \temp_ALUop_output~0_combout ;
wire \temp_ALUop_output~1_combout ;
wire \temp_ALUsrc_output~0_combout ;
wire \temp_ALUop_output~3_combout ;
wire \temp_imemload_output~0_combout ;
wire \temp_imemload_output~1_combout ;
wire \temp_ALUsrc_output~1_combout ;
wire \temp_ALUsrc_output[0]~2_combout ;
wire \temp_branch_output~1_combout ;
wire \temp_ALUsrc_output~4_combout ;
wire \temp_rdat_two_output~0_combout ;
wire \temp_imemload_output~2_combout ;
wire \temp_imemload_output~3_combout ;
wire \temp_imemload_output~4_combout ;
wire \temp_imemload_output~5_combout ;
wire \temp_imemload_output~6_combout ;
wire \temp_imemload_output~7_combout ;
wire \temp_imemload_output~8_combout ;
wire \temp_imemload_output~9_combout ;
wire \temp_imemload_output~10_combout ;
wire \temp_imemload_output~11_combout ;
wire \temp_rdat_one_output~0_combout ;
wire \temp_ALUop_output~4_combout ;
wire \temp_ALUop_output~5_combout ;
wire \temp_ALUop_output~6_combout ;
wire \temp_imemload_output~12_combout ;
wire \temp_imemload_output~13_combout ;
wire \temp_rdat_two_output~1_combout ;
wire \temp_rdat_one_output~1_combout ;
wire \temp_rdat_one_output~2_combout ;
wire \temp_rdat_one_output~3_combout ;
wire \temp_rdat_one_output~4_combout ;
wire \temp_imemload_output~14_combout ;
wire \temp_imemload_output~15_combout ;
wire \temp_rdat_two_output~2_combout ;
wire \temp_rdat_one_output~5_combout ;
wire \temp_rdat_one_output~6_combout ;
wire \temp_rdat_one_output~7_combout ;
wire \temp_rdat_one_output~8_combout ;
wire \temp_imemload_output~16_combout ;
wire \temp_imemload_output~17_combout ;
wire \temp_rdat_two_output~3_combout ;
wire \temp_rdat_one_output~9_combout ;
wire \temp_rdat_one_output~10_combout ;
wire \temp_rdat_one_output~11_combout ;
wire \temp_rdat_one_output~12_combout ;
wire \temp_rdat_one_output~13_combout ;
wire \temp_rdat_one_output~14_combout ;
wire \temp_rdat_one_output~15_combout ;
wire \temp_rdat_one_output~16_combout ;
wire \temp_imemload_output~18_combout ;
wire \temp_imemload_output~19_combout ;
wire \temp_rdat_two_output~4_combout ;
wire \temp_rdat_one_output~17_combout ;
wire \temp_rdat_one_output~18_combout ;
wire \temp_rdat_one_output~19_combout ;
wire \temp_rdat_one_output~20_combout ;
wire \temp_rdat_one_output~21_combout ;
wire \temp_rdat_one_output~22_combout ;
wire \temp_rdat_one_output~23_combout ;
wire \temp_rdat_one_output~24_combout ;
wire \temp_rdat_one_output~25_combout ;
wire \temp_rdat_one_output~26_combout ;
wire \temp_rdat_one_output~27_combout ;
wire \temp_rdat_one_output~28_combout ;
wire \temp_rdat_one_output~29_combout ;
wire \temp_rdat_one_output~30_combout ;
wire \temp_rdat_one_output~31_combout ;
wire \temp_rdat_two_output~5_combout ;
wire \temp_imemload_output~20_combout ;
wire \temp_rdat_two_output~6_combout ;
wire \temp_imemload_output~21_combout ;
wire \temp_rdat_two_output~7_combout ;
wire \temp_rdat_two_output~8_combout ;
wire \temp_rdat_two_output~9_combout ;
wire \temp_rdat_two_output~10_combout ;
wire \temp_rdat_two_output~11_combout ;
wire \temp_rdat_two_output~12_combout ;
wire \temp_rdat_two_output~13_combout ;
wire \temp_rdat_two_output~14_combout ;
wire \temp_rdat_two_output~15_combout ;
wire \temp_rdat_two_output~16_combout ;
wire \temp_rdat_two_output~17_combout ;
wire \temp_rdat_two_output~18_combout ;
wire \temp_rdat_two_output~19_combout ;
wire \temp_rdat_two_output~20_combout ;
wire \temp_rdat_two_output~21_combout ;
wire \temp_rdat_two_output~22_combout ;
wire \temp_imemload_output~22_combout ;
wire \temp_rdat_two_output~23_combout ;
wire \temp_rdat_two_output~24_combout ;
wire \temp_rdat_two_output~25_combout ;
wire \temp_rdat_two_output~26_combout ;
wire \temp_rdat_two_output~27_combout ;
wire \temp_rdat_two_output~28_combout ;
wire \temp_rdat_two_output~29_combout ;
wire \temp_imemload_output~23_combout ;
wire \temp_rdat_two_output~30_combout ;
wire \temp_imemload_output~24_combout ;
wire \temp_rdat_two_output~31_combout ;
wire \temp_imemload_output~25_combout ;
wire \temp_ALUop_output~7_combout ;
wire \temp_ALUop_output~8_combout ;
wire \temp_ALUop_output~9_combout ;
wire \temp_ALUop_output~10_combout ;
wire \temp_ALUop_output~11_combout ;
wire \temp_request_dmemREN_output~0_combout ;
wire \temp_request_dmemREN_output~1_combout ;
wire \temp_request_dmemWEN_output~0_combout ;
wire \temp_regdst_output~0_combout ;
wire \temp_regwrite_output~0_combout ;
wire \temp_regwrite_output~1_combout ;
wire \temp_regdst_output~1_combout ;
wire \temp_regdst_output~2_combout ;
wire \temp_request_dmemREN_output~2_combout ;
wire \temp_memtoreg_output~0_combout ;
wire \temp_imemload_output~26_combout ;
wire \temp_imemload_output~27_combout ;
wire \temp_imemload_output~28_combout ;
wire \temp_imemload_output~29_combout ;
wire \temp_imemload_output~30_combout ;
wire \temp_imemload_output~31_combout ;
wire \temp_branch_output~2_combout ;
wire \temp_branch_output~3_combout ;
wire \temp_NPC_output~0_combout ;
wire \temp_pcselect_output~0_combout ;
wire \temp_pcselect_output~1_combout ;
wire \temp_pcselect_output~2_combout ;
wire \temp_pcselect_output~3_combout ;
wire \temp_NPC_output~1_combout ;
wire \temp_NPC_output~2_combout ;
wire \temp_NPC_output~3_combout ;
wire \temp_NPC_output~4_combout ;
wire \temp_NPC_output~5_combout ;
wire \temp_NPC_output~6_combout ;
wire \temp_NPC_output~7_combout ;
wire \temp_NPC_output~8_combout ;
wire \temp_NPC_output~9_combout ;
wire \temp_NPC_output~10_combout ;
wire \temp_NPC_output~11_combout ;
wire \temp_NPC_output~12_combout ;
wire \temp_NPC_output~13_combout ;
wire \temp_NPC_output~14_combout ;
wire \temp_NPC_output~15_combout ;
wire \temp_NPC_output~16_combout ;
wire \temp_NPC_output~17_combout ;
wire \temp_NPC_output~18_combout ;
wire \temp_NPC_output~19_combout ;
wire \temp_NPC_output~20_combout ;
wire \temp_NPC_output~21_combout ;
wire \temp_NPC_output[21]~feeder_combout ;
wire \temp_NPC_output~22_combout ;
wire \temp_NPC_output~23_combout ;
wire \temp_NPC_output~24_combout ;
wire \temp_NPC_output~25_combout ;
wire \temp_NPC_output~26_combout ;
wire \temp_NPC_output~27_combout ;
wire \temp_NPC_output~28_combout ;
wire \temp_NPC_output~29_combout ;
wire \temp_NPC_output~30_combout ;
wire \temp_NPC_output~31_combout ;


// Location: FF_X66_Y36_N21
dffeas \temp_signzerovalue_output[16] (
	.clk(CLK),
	.d(extended_imm_161),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(id_ex_flush),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_signzerovalue_output_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_signzerovalue_output[16] .is_wysiwyg = "true";
defparam \temp_signzerovalue_output[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N13
dffeas temp_halt_out_output(
	.clk(CLK),
	.d(halt_out1),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(id_ex_flush),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_halt_out_output1),
	.prn(vcc));
// synopsys translate_off
defparam temp_halt_out_output.is_wysiwyg = "true";
defparam temp_halt_out_output.power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N31
dffeas \temp_ALUop_output[0] (
	.clk(CLK),
	.d(\temp_ALUop_output~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_ALUop_output_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_ALUop_output[0] .is_wysiwyg = "true";
defparam \temp_ALUop_output[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N21
dffeas \temp_imemload_output[1] (
	.clk(CLK),
	.d(\temp_imemload_output~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[1] .is_wysiwyg = "true";
defparam \temp_imemload_output[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N21
dffeas \temp_imemload_output[7] (
	.clk(CLK),
	.d(\temp_imemload_output~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[7] .is_wysiwyg = "true";
defparam \temp_imemload_output[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N15
dffeas \temp_ALUsrc_output[1] (
	.clk(CLK),
	.d(\temp_ALUsrc_output~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_ALUsrc_output_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_ALUsrc_output[1] .is_wysiwyg = "true";
defparam \temp_ALUsrc_output[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y36_N17
dffeas \temp_ALUsrc_output[0] (
	.clk(CLK),
	.d(\temp_ALUsrc_output~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_ALUsrc_output_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_ALUsrc_output[0] .is_wysiwyg = "true";
defparam \temp_ALUsrc_output[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N1
dffeas \temp_rdat_two_output[1] (
	.clk(CLK),
	.d(\temp_rdat_two_output~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[1] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y44_N17
dffeas \temp_imemload_output[17] (
	.clk(CLK),
	.d(\temp_imemload_output~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[17] .is_wysiwyg = "true";
defparam \temp_imemload_output[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y44_N19
dffeas \temp_imemload_output[16] (
	.clk(CLK),
	.d(\temp_imemload_output~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[16] .is_wysiwyg = "true";
defparam \temp_imemload_output[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y44_N27
dffeas \temp_imemload_output[18] (
	.clk(CLK),
	.d(\temp_imemload_output~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[18] .is_wysiwyg = "true";
defparam \temp_imemload_output[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y44_N17
dffeas \temp_imemload_output[19] (
	.clk(CLK),
	.d(\temp_imemload_output~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[19] .is_wysiwyg = "true";
defparam \temp_imemload_output[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N17
dffeas \temp_imemload_output[20] (
	.clk(CLK),
	.d(\temp_imemload_output~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[20] .is_wysiwyg = "true";
defparam \temp_imemload_output[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y44_N5
dffeas \temp_imemload_output[22] (
	.clk(CLK),
	.d(\temp_imemload_output~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[22] .is_wysiwyg = "true";
defparam \temp_imemload_output[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y44_N27
dffeas \temp_imemload_output[21] (
	.clk(CLK),
	.d(\temp_imemload_output~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[21] .is_wysiwyg = "true";
defparam \temp_imemload_output[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N3
dffeas \temp_imemload_output[23] (
	.clk(CLK),
	.d(\temp_imemload_output~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[23] .is_wysiwyg = "true";
defparam \temp_imemload_output[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N5
dffeas \temp_imemload_output[24] (
	.clk(CLK),
	.d(\temp_imemload_output~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[24] .is_wysiwyg = "true";
defparam \temp_imemload_output[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N17
dffeas \temp_imemload_output[25] (
	.clk(CLK),
	.d(\temp_imemload_output~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[25] .is_wysiwyg = "true";
defparam \temp_imemload_output[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y44_N27
dffeas \temp_rdat_one_output[1] (
	.clk(CLK),
	.d(\temp_rdat_one_output~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[1] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N17
dffeas \temp_ALUop_output[1] (
	.clk(CLK),
	.d(\temp_ALUop_output~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_ALUop_output_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_ALUop_output[1] .is_wysiwyg = "true";
defparam \temp_ALUop_output[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N5
dffeas \temp_imemload_output[0] (
	.clk(CLK),
	.d(\temp_imemload_output~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[0] .is_wysiwyg = "true";
defparam \temp_imemload_output[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N27
dffeas \temp_imemload_output[6] (
	.clk(CLK),
	.d(\temp_imemload_output~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[6] .is_wysiwyg = "true";
defparam \temp_imemload_output[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N5
dffeas \temp_rdat_two_output[0] (
	.clk(CLK),
	.d(\temp_rdat_two_output~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[0] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N29
dffeas \temp_rdat_one_output[0] (
	.clk(CLK),
	.d(\temp_rdat_one_output~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[0] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y42_N31
dffeas \temp_rdat_one_output[2] (
	.clk(CLK),
	.d(\temp_rdat_one_output~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[2] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N1
dffeas \temp_rdat_one_output[4] (
	.clk(CLK),
	.d(\temp_rdat_one_output~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[4] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N19
dffeas \temp_rdat_one_output[3] (
	.clk(CLK),
	.d(\temp_rdat_one_output~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[3] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y44_N29
dffeas \temp_imemload_output[2] (
	.clk(CLK),
	.d(\temp_imemload_output~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[2] .is_wysiwyg = "true";
defparam \temp_imemload_output[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N17
dffeas \temp_imemload_output[8] (
	.clk(CLK),
	.d(\temp_imemload_output~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[8] .is_wysiwyg = "true";
defparam \temp_imemload_output[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N29
dffeas \temp_rdat_two_output[2] (
	.clk(CLK),
	.d(\temp_rdat_two_output~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[2] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N9
dffeas \temp_rdat_one_output[8] (
	.clk(CLK),
	.d(\temp_rdat_one_output~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[8] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N25
dffeas \temp_rdat_one_output[7] (
	.clk(CLK),
	.d(\temp_rdat_one_output~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[7] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y42_N27
dffeas \temp_rdat_one_output[6] (
	.clk(CLK),
	.d(\temp_rdat_one_output~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[6] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N15
dffeas \temp_rdat_one_output[5] (
	.clk(CLK),
	.d(\temp_rdat_one_output~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[5] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N27
dffeas \temp_imemload_output[3] (
	.clk(CLK),
	.d(\temp_imemload_output~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[3] .is_wysiwyg = "true";
defparam \temp_imemload_output[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N9
dffeas \temp_imemload_output[9] (
	.clk(CLK),
	.d(\temp_imemload_output~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[9] .is_wysiwyg = "true";
defparam \temp_imemload_output[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N17
dffeas \temp_rdat_two_output[3] (
	.clk(CLK),
	.d(\temp_rdat_two_output~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[3] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N1
dffeas \temp_rdat_one_output[16] (
	.clk(CLK),
	.d(\temp_rdat_one_output~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[16] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N25
dffeas \temp_rdat_one_output[14] (
	.clk(CLK),
	.d(\temp_rdat_one_output~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[14] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N23
dffeas \temp_rdat_one_output[15] (
	.clk(CLK),
	.d(\temp_rdat_one_output~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[15] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N31
dffeas \temp_rdat_one_output[13] (
	.clk(CLK),
	.d(\temp_rdat_one_output~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[13] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y43_N25
dffeas \temp_rdat_one_output[12] (
	.clk(CLK),
	.d(\temp_rdat_one_output~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[12] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N31
dffeas \temp_rdat_one_output[10] (
	.clk(CLK),
	.d(\temp_rdat_one_output~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[10] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N15
dffeas \temp_rdat_one_output[11] (
	.clk(CLK),
	.d(\temp_rdat_one_output~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[11] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N19
dffeas \temp_rdat_one_output[9] (
	.clk(CLK),
	.d(\temp_rdat_one_output~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[9] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N29
dffeas \temp_imemload_output[4] (
	.clk(CLK),
	.d(\temp_imemload_output~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[4] .is_wysiwyg = "true";
defparam \temp_imemload_output[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N23
dffeas \temp_imemload_output[10] (
	.clk(CLK),
	.d(\temp_imemload_output~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[10] .is_wysiwyg = "true";
defparam \temp_imemload_output[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N17
dffeas \temp_rdat_two_output[4] (
	.clk(CLK),
	.d(\temp_rdat_two_output~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[4] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N3
dffeas \temp_rdat_one_output[31] (
	.clk(CLK),
	.d(\temp_rdat_one_output~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[31] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N3
dffeas \temp_rdat_one_output[30] (
	.clk(CLK),
	.d(\temp_rdat_one_output~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[30] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N1
dffeas \temp_rdat_one_output[29] (
	.clk(CLK),
	.d(\temp_rdat_one_output~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[29] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N29
dffeas \temp_rdat_one_output[26] (
	.clk(CLK),
	.d(\temp_rdat_one_output~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[26] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N1
dffeas \temp_rdat_one_output[25] (
	.clk(CLK),
	.d(\temp_rdat_one_output~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[25] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N13
dffeas \temp_rdat_one_output[28] (
	.clk(CLK),
	.d(\temp_rdat_one_output~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[28] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N1
dffeas \temp_rdat_one_output[27] (
	.clk(CLK),
	.d(\temp_rdat_one_output~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[27] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N9
dffeas \temp_rdat_one_output[17] (
	.clk(CLK),
	.d(\temp_rdat_one_output~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[17] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N11
dffeas \temp_rdat_one_output[20] (
	.clk(CLK),
	.d(\temp_rdat_one_output~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[20] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N11
dffeas \temp_rdat_one_output[19] (
	.clk(CLK),
	.d(\temp_rdat_one_output~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[19] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N15
dffeas \temp_rdat_one_output[18] (
	.clk(CLK),
	.d(\temp_rdat_one_output~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[18] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N15
dffeas \temp_rdat_one_output[24] (
	.clk(CLK),
	.d(\temp_rdat_one_output~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[24] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N17
dffeas \temp_rdat_one_output[23] (
	.clk(CLK),
	.d(\temp_rdat_one_output~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[23] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N25
dffeas \temp_rdat_one_output[22] (
	.clk(CLK),
	.d(\temp_rdat_one_output~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[22] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N15
dffeas \temp_rdat_one_output[21] (
	.clk(CLK),
	.d(\temp_rdat_one_output~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_one_output_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_one_output[21] .is_wysiwyg = "true";
defparam \temp_rdat_one_output[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N19
dffeas \temp_rdat_two_output[15] (
	.clk(CLK),
	.d(\temp_rdat_two_output~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[15] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N7
dffeas \temp_imemload_output[15] (
	.clk(CLK),
	.d(\temp_imemload_output~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[15] .is_wysiwyg = "true";
defparam \temp_imemload_output[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N5
dffeas \temp_rdat_two_output[12] (
	.clk(CLK),
	.d(\temp_rdat_two_output~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[12] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N27
dffeas \temp_imemload_output[12] (
	.clk(CLK),
	.d(\temp_imemload_output~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[12] .is_wysiwyg = "true";
defparam \temp_imemload_output[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N13
dffeas \temp_rdat_two_output[27] (
	.clk(CLK),
	.d(\temp_rdat_two_output~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[27] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N5
dffeas \temp_rdat_two_output[18] (
	.clk(CLK),
	.d(\temp_rdat_two_output~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[18] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N23
dffeas \temp_rdat_two_output[17] (
	.clk(CLK),
	.d(\temp_rdat_two_output~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[17] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N3
dffeas \temp_rdat_two_output[16] (
	.clk(CLK),
	.d(\temp_rdat_two_output~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[16] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N23
dffeas \temp_rdat_two_output[31] (
	.clk(CLK),
	.d(\temp_rdat_two_output~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[31] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N31
dffeas \temp_rdat_two_output[30] (
	.clk(CLK),
	.d(\temp_rdat_two_output~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[30] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N13
dffeas \temp_rdat_two_output[29] (
	.clk(CLK),
	.d(\temp_rdat_two_output~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[29] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N5
dffeas \temp_rdat_two_output[28] (
	.clk(CLK),
	.d(\temp_rdat_two_output~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[28] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N25
dffeas \temp_rdat_two_output[26] (
	.clk(CLK),
	.d(\temp_rdat_two_output~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[26] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N15
dffeas \temp_rdat_two_output[25] (
	.clk(CLK),
	.d(\temp_rdat_two_output~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[25] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N29
dffeas \temp_rdat_two_output[24] (
	.clk(CLK),
	.d(\temp_rdat_two_output~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[24] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N5
dffeas \temp_rdat_two_output[23] (
	.clk(CLK),
	.d(\temp_rdat_two_output~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[23] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N3
dffeas \temp_rdat_two_output[22] (
	.clk(CLK),
	.d(\temp_rdat_two_output~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[22] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N25
dffeas \temp_rdat_two_output[21] (
	.clk(CLK),
	.d(\temp_rdat_two_output~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[21] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N17
dffeas \temp_rdat_two_output[20] (
	.clk(CLK),
	.d(\temp_rdat_two_output~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[20] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N29
dffeas \temp_rdat_two_output[19] (
	.clk(CLK),
	.d(\temp_rdat_two_output~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[19] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N21
dffeas \temp_imemload_output[14] (
	.clk(CLK),
	.d(\temp_imemload_output~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[14] .is_wysiwyg = "true";
defparam \temp_imemload_output[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N21
dffeas \temp_rdat_two_output[10] (
	.clk(CLK),
	.d(\temp_rdat_two_output~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[10] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N13
dffeas \temp_rdat_two_output[14] (
	.clk(CLK),
	.d(\temp_rdat_two_output~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[14] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N13
dffeas \temp_rdat_two_output[9] (
	.clk(CLK),
	.d(\temp_rdat_two_output~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[9] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N7
dffeas \temp_rdat_two_output[8] (
	.clk(CLK),
	.d(\temp_rdat_two_output~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[8] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N19
dffeas \temp_rdat_two_output[7] (
	.clk(CLK),
	.d(\temp_rdat_two_output~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[7] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y42_N17
dffeas \temp_rdat_two_output[6] (
	.clk(CLK),
	.d(\temp_rdat_two_output~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[6] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N21
dffeas \temp_rdat_two_output[5] (
	.clk(CLK),
	.d(\temp_rdat_two_output~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[5] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N31
dffeas \temp_imemload_output[5] (
	.clk(CLK),
	.d(\temp_imemload_output~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[5] .is_wysiwyg = "true";
defparam \temp_imemload_output[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N11
dffeas \temp_rdat_two_output[13] (
	.clk(CLK),
	.d(\temp_rdat_two_output~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[13] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N21
dffeas \temp_imemload_output[13] (
	.clk(CLK),
	.d(\temp_imemload_output~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[13] .is_wysiwyg = "true";
defparam \temp_imemload_output[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N31
dffeas \temp_rdat_two_output[11] (
	.clk(CLK),
	.d(\temp_rdat_two_output~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_rdat_two_output_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_rdat_two_output[11] .is_wysiwyg = "true";
defparam \temp_rdat_two_output[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N25
dffeas \temp_imemload_output[11] (
	.clk(CLK),
	.d(\temp_imemload_output~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[11] .is_wysiwyg = "true";
defparam \temp_imemload_output[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N11
dffeas \temp_ALUop_output[2] (
	.clk(CLK),
	.d(\temp_ALUop_output~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_ALUop_output_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_ALUop_output[2] .is_wysiwyg = "true";
defparam \temp_ALUop_output[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N29
dffeas \temp_ALUop_output[3] (
	.clk(CLK),
	.d(\temp_ALUop_output~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_ALUop_output_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_ALUop_output[3] .is_wysiwyg = "true";
defparam \temp_ALUop_output[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y44_N21
dffeas temp_request_dmemREN_output(
	.clk(CLK),
	.d(\temp_request_dmemREN_output~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_request_dmemREN_output1),
	.prn(vcc));
// synopsys translate_off
defparam temp_request_dmemREN_output.is_wysiwyg = "true";
defparam temp_request_dmemREN_output.power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y36_N19
dffeas temp_request_dmemWEN_output(
	.clk(CLK),
	.d(\temp_request_dmemWEN_output~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_request_dmemWEN_output1),
	.prn(vcc));
// synopsys translate_off
defparam temp_request_dmemWEN_output.is_wysiwyg = "true";
defparam temp_request_dmemWEN_output.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N22
cycloneive_lcell_comb \temp_branch_output~0 (
// Equation(s):
// temp_branch_output1 = (!temp_imemload_output_26 & !temp_imemload_output_27)

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_imemload_output_26),
	.datad(temp_imemload_output_27),
	.cin(gnd),
	.combout(temp_branch_output1),
	.cout());
// synopsys translate_off
defparam \temp_branch_output~0 .lut_mask = 16'h000F;
defparam \temp_branch_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N28
cycloneive_lcell_comb \temp_ALUsrc_output~3 (
// Equation(s):
// temp_ALUsrc_output = (temp_imemload_output_27 & (temp_imemload_output_31 & (temp_imemload_output_26 & !temp_imemload_output_28)))

	.dataa(temp_imemload_output_27),
	.datab(temp_imemload_output_31),
	.datac(temp_imemload_output_26),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(temp_ALUsrc_output),
	.cout());
// synopsys translate_off
defparam \temp_ALUsrc_output~3 .lut_mask = 16'h0080;
defparam \temp_ALUsrc_output~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y36_N1
dffeas temp_regwrite_output(
	.clk(CLK),
	.d(\temp_regwrite_output~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_regwrite_output1),
	.prn(vcc));
// synopsys translate_off
defparam temp_regwrite_output.is_wysiwyg = "true";
defparam temp_regwrite_output.power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y44_N29
dffeas \temp_regdst_output[1] (
	.clk(CLK),
	.d(\temp_regdst_output~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_regdst_output_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_regdst_output[1] .is_wysiwyg = "true";
defparam \temp_regdst_output[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N11
dffeas \temp_regdst_output[0] (
	.clk(CLK),
	.d(\temp_regdst_output~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_regdst_output_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_regdst_output[0] .is_wysiwyg = "true";
defparam \temp_regdst_output[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y44_N11
dffeas \temp_memtoreg_output[0] (
	.clk(CLK),
	.d(\temp_request_dmemREN_output~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_memtoreg_output_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_memtoreg_output[0] .is_wysiwyg = "true";
defparam \temp_memtoreg_output[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N27
dffeas \temp_memtoreg_output[1] (
	.clk(CLK),
	.d(\temp_memtoreg_output~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_memtoreg_output_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_memtoreg_output[1] .is_wysiwyg = "true";
defparam \temp_memtoreg_output[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N11
dffeas \temp_imemload_output[31] (
	.clk(CLK),
	.d(\temp_imemload_output~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_311),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[31] .is_wysiwyg = "true";
defparam \temp_imemload_output[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N3
dffeas \temp_imemload_output[30] (
	.clk(CLK),
	.d(\temp_imemload_output~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_301),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[30] .is_wysiwyg = "true";
defparam \temp_imemload_output[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N21
dffeas \temp_imemload_output[29] (
	.clk(CLK),
	.d(\temp_imemload_output~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_291),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[29] .is_wysiwyg = "true";
defparam \temp_imemload_output[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y42_N25
dffeas \temp_imemload_output[27] (
	.clk(CLK),
	.d(\temp_imemload_output~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_271),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[27] .is_wysiwyg = "true";
defparam \temp_imemload_output[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y42_N11
dffeas \temp_imemload_output[26] (
	.clk(CLK),
	.d(\temp_imemload_output~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_261),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[26] .is_wysiwyg = "true";
defparam \temp_imemload_output[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y42_N5
dffeas \temp_imemload_output[28] (
	.clk(CLK),
	.d(\temp_imemload_output~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_281),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[28] .is_wysiwyg = "true";
defparam \temp_imemload_output[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N19
dffeas temp_branch_output(
	.clk(CLK),
	.d(\temp_branch_output~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branch_output2),
	.prn(vcc));
// synopsys translate_off
defparam temp_branch_output.is_wysiwyg = "true";
defparam temp_branch_output.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N3
dffeas \temp_NPC_output[1] (
	.clk(CLK),
	.d(\temp_NPC_output~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[1] .is_wysiwyg = "true";
defparam \temp_NPC_output[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N9
dffeas \temp_pcselect_output[1] (
	.clk(CLK),
	.d(\temp_pcselect_output~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_pcselect_output_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_pcselect_output[1] .is_wysiwyg = "true";
defparam \temp_pcselect_output[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N25
dffeas \temp_pcselect_output[0] (
	.clk(CLK),
	.d(\temp_pcselect_output~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_pcselect_output_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_pcselect_output[0] .is_wysiwyg = "true";
defparam \temp_pcselect_output[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N25
dffeas \temp_NPC_output[0] (
	.clk(CLK),
	.d(\temp_NPC_output~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[0] .is_wysiwyg = "true";
defparam \temp_NPC_output[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N11
dffeas \temp_NPC_output[2] (
	.clk(CLK),
	.d(\temp_NPC_output~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[2] .is_wysiwyg = "true";
defparam \temp_NPC_output[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N29
dffeas \temp_NPC_output[3] (
	.clk(CLK),
	.d(\temp_NPC_output~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[3] .is_wysiwyg = "true";
defparam \temp_NPC_output[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N25
dffeas \temp_NPC_output[5] (
	.clk(CLK),
	.d(\temp_NPC_output~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[5] .is_wysiwyg = "true";
defparam \temp_NPC_output[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y44_N21
dffeas \temp_NPC_output[4] (
	.clk(CLK),
	.d(\temp_NPC_output~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[4] .is_wysiwyg = "true";
defparam \temp_NPC_output[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N13
dffeas \temp_NPC_output[7] (
	.clk(CLK),
	.d(\temp_NPC_output~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[7] .is_wysiwyg = "true";
defparam \temp_NPC_output[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N11
dffeas \temp_NPC_output[6] (
	.clk(CLK),
	.d(\temp_NPC_output~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[6] .is_wysiwyg = "true";
defparam \temp_NPC_output[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N29
dffeas \temp_NPC_output[9] (
	.clk(CLK),
	.d(\temp_NPC_output~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[9] .is_wysiwyg = "true";
defparam \temp_NPC_output[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N7
dffeas \temp_NPC_output[8] (
	.clk(CLK),
	.d(\temp_NPC_output~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[8] .is_wysiwyg = "true";
defparam \temp_NPC_output[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N3
dffeas \temp_NPC_output[11] (
	.clk(CLK),
	.d(\temp_NPC_output~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[11] .is_wysiwyg = "true";
defparam \temp_NPC_output[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N21
dffeas \temp_NPC_output[10] (
	.clk(CLK),
	.d(\temp_NPC_output~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[10] .is_wysiwyg = "true";
defparam \temp_NPC_output[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N17
dffeas \temp_NPC_output[13] (
	.clk(CLK),
	.d(\temp_NPC_output~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[13] .is_wysiwyg = "true";
defparam \temp_NPC_output[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N15
dffeas \temp_NPC_output[12] (
	.clk(CLK),
	.d(\temp_NPC_output~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[12] .is_wysiwyg = "true";
defparam \temp_NPC_output[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N11
dffeas \temp_NPC_output[15] (
	.clk(CLK),
	.d(\temp_NPC_output~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[15] .is_wysiwyg = "true";
defparam \temp_NPC_output[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N17
dffeas \temp_NPC_output[14] (
	.clk(CLK),
	.d(\temp_NPC_output~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[14] .is_wysiwyg = "true";
defparam \temp_NPC_output[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N1
dffeas \temp_NPC_output[17] (
	.clk(CLK),
	.d(\temp_NPC_output~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[17] .is_wysiwyg = "true";
defparam \temp_NPC_output[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N1
dffeas \temp_NPC_output[16] (
	.clk(CLK),
	.d(\temp_NPC_output~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[16] .is_wysiwyg = "true";
defparam \temp_NPC_output[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N13
dffeas \temp_NPC_output[19] (
	.clk(CLK),
	.d(\temp_NPC_output~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[19] .is_wysiwyg = "true";
defparam \temp_NPC_output[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N19
dffeas \temp_NPC_output[18] (
	.clk(CLK),
	.d(\temp_NPC_output~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[18] .is_wysiwyg = "true";
defparam \temp_NPC_output[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N19
dffeas \temp_NPC_output[20] (
	.clk(CLK),
	.d(\temp_NPC_output~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[20] .is_wysiwyg = "true";
defparam \temp_NPC_output[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N15
dffeas \temp_NPC_output[21] (
	.clk(CLK),
	.d(\temp_NPC_output[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[21] .is_wysiwyg = "true";
defparam \temp_NPC_output[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N31
dffeas \temp_NPC_output[23] (
	.clk(CLK),
	.d(\temp_NPC_output~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[23] .is_wysiwyg = "true";
defparam \temp_NPC_output[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y44_N15
dffeas \temp_NPC_output[22] (
	.clk(CLK),
	.d(\temp_NPC_output~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[22] .is_wysiwyg = "true";
defparam \temp_NPC_output[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N1
dffeas \temp_NPC_output[25] (
	.clk(CLK),
	.d(\temp_NPC_output~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[25] .is_wysiwyg = "true";
defparam \temp_NPC_output[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y44_N21
dffeas \temp_NPC_output[24] (
	.clk(CLK),
	.d(\temp_NPC_output~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[24] .is_wysiwyg = "true";
defparam \temp_NPC_output[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N1
dffeas \temp_NPC_output[26] (
	.clk(CLK),
	.d(\temp_NPC_output~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[26] .is_wysiwyg = "true";
defparam \temp_NPC_output[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N21
dffeas \temp_NPC_output[27] (
	.clk(CLK),
	.d(\temp_NPC_output~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[27] .is_wysiwyg = "true";
defparam \temp_NPC_output[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N17
dffeas \temp_NPC_output[29] (
	.clk(CLK),
	.d(\temp_NPC_output~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[29] .is_wysiwyg = "true";
defparam \temp_NPC_output[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N15
dffeas \temp_NPC_output[28] (
	.clk(CLK),
	.d(\temp_NPC_output~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[28] .is_wysiwyg = "true";
defparam \temp_NPC_output[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N31
dffeas \temp_NPC_output[31] (
	.clk(CLK),
	.d(\temp_NPC_output~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[31] .is_wysiwyg = "true";
defparam \temp_NPC_output[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N25
dffeas \temp_NPC_output[30] (
	.clk(CLK),
	.d(\temp_NPC_output~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[30] .is_wysiwyg = "true";
defparam \temp_NPC_output[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N12
cycloneive_lcell_comb \temp_ALUop_output~2 (
// Equation(s):
// \temp_ALUop_output~2_combout  = (Equal31 & ((temp_imemload_output_1) # ((temp_imemload_output_5 & WideOr2)))) # (!Equal31 & (temp_imemload_output_5 & (WideOr2)))

	.dataa(Equal31),
	.datab(temp_imemload_output_51),
	.datac(WideOr2),
	.datad(temp_imemload_output_110),
	.cin(gnd),
	.combout(\temp_ALUop_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~2 .lut_mask = 16'hEAC0;
defparam \temp_ALUop_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N16
cycloneive_lcell_comb \temp_ALUop_output~0 (
// Equation(s):
// \temp_ALUop_output~0_combout  = (!ex_mem_flush3 & (!use_after_load & !Equal32))

	.dataa(ex_mem_flush),
	.datab(use_after_load),
	.datac(gnd),
	.datad(Equal32),
	.cin(gnd),
	.combout(\temp_ALUop_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~0 .lut_mask = 16'h0011;
defparam \temp_ALUop_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N26
cycloneive_lcell_comb \temp_ALUop_output~1 (
// Equation(s):
// \temp_ALUop_output~1_combout  = (extended_imm_16 & (WideOr8 & !temp_imemload_output_31))

	.dataa(extended_imm_16),
	.datab(WideOr8),
	.datac(temp_imemload_output_31),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_ALUop_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~1 .lut_mask = 16'h0808;
defparam \temp_ALUop_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N4
cycloneive_lcell_comb \temp_ALUsrc_output~0 (
// Equation(s):
// \temp_ALUsrc_output~0_combout  = (temp_branch_output1 & (Equal3 & (!temp_imemload_output_4 & !Equal32)))

	.dataa(temp_branch_output1),
	.datab(Equal3),
	.datac(temp_imemload_output_41),
	.datad(Equal32),
	.cin(gnd),
	.combout(\temp_ALUsrc_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUsrc_output~0 .lut_mask = 16'h0008;
defparam \temp_ALUsrc_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N30
cycloneive_lcell_comb \temp_ALUop_output~3 (
// Equation(s):
// \temp_ALUop_output~3_combout  = (\temp_ALUop_output~0_combout  & ((\temp_ALUop_output~1_combout ) # ((\temp_ALUop_output~2_combout  & \temp_ALUsrc_output~0_combout ))))

	.dataa(\temp_ALUop_output~2_combout ),
	.datab(\temp_ALUop_output~0_combout ),
	.datac(\temp_ALUop_output~1_combout ),
	.datad(\temp_ALUsrc_output~0_combout ),
	.cin(gnd),
	.combout(\temp_ALUop_output~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~3 .lut_mask = 16'hC8C0;
defparam \temp_ALUop_output~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N20
cycloneive_lcell_comb \temp_imemload_output~0 (
// Equation(s):
// \temp_imemload_output~0_combout  = (!use_after_load & (temp_imemload_output_1 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(use_after_load),
	.datac(temp_imemload_output_110),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_imemload_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~0 .lut_mask = 16'h0030;
defparam \temp_imemload_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N20
cycloneive_lcell_comb \temp_imemload_output~1 (
// Equation(s):
// \temp_imemload_output~1_combout  = (!ex_mem_flush3 & (!use_after_load & temp_imemload_output_7))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(use_after_load),
	.datad(temp_imemload_output_71),
	.cin(gnd),
	.combout(\temp_imemload_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~1 .lut_mask = 16'h0500;
defparam \temp_imemload_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N14
cycloneive_lcell_comb \temp_ALUsrc_output~1 (
// Equation(s):
// \temp_ALUsrc_output~1_combout  = (Equal31 & (\temp_ALUsrc_output~0_combout  & !id_ex_flush1))

	.dataa(Equal31),
	.datab(\temp_ALUsrc_output~0_combout ),
	.datac(gnd),
	.datad(id_ex_flush),
	.cin(gnd),
	.combout(\temp_ALUsrc_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUsrc_output~1 .lut_mask = 16'h0088;
defparam \temp_ALUsrc_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N18
cycloneive_lcell_comb \temp_ALUsrc_output[0]~2 (
// Equation(s):
// \temp_ALUsrc_output[0]~2_combout  = (id_ex_flush1) # ((Equal32) # ((temp_branch_output1 & Equal3)))

	.dataa(temp_branch_output1),
	.datab(id_ex_flush),
	.datac(Equal3),
	.datad(Equal32),
	.cin(gnd),
	.combout(\temp_ALUsrc_output[0]~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUsrc_output[0]~2 .lut_mask = 16'hFFEC;
defparam \temp_ALUsrc_output[0]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N28
cycloneive_lcell_comb \temp_branch_output~1 (
// Equation(s):
// \temp_branch_output~1_combout  = (!temp_imemload_output_30 & !\temp_ALUsrc_output[0]~2_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_imemload_output_30),
	.datad(\temp_ALUsrc_output[0]~2_combout ),
	.cin(gnd),
	.combout(\temp_branch_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_branch_output~1 .lut_mask = 16'h000F;
defparam \temp_branch_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N16
cycloneive_lcell_comb \temp_ALUsrc_output~4 (
// Equation(s):
// \temp_ALUsrc_output~4_combout  = (\temp_branch_output~1_combout  & ((temp_imemload_output_29 & ((WideOr4))) # (!temp_imemload_output_29 & (temp_ALUsrc_output))))

	.dataa(temp_ALUsrc_output),
	.datab(\temp_branch_output~1_combout ),
	.datac(temp_imemload_output_29),
	.datad(WideOr4),
	.cin(gnd),
	.combout(\temp_ALUsrc_output~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUsrc_output~4 .lut_mask = 16'hC808;
defparam \temp_ALUsrc_output~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N0
cycloneive_lcell_comb \temp_rdat_two_output~0 (
// Equation(s):
// \temp_rdat_two_output~0_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux62)) # (!temp_imemload_output_20 & ((Mux621)))))

	.dataa(id_ex_flush),
	.datab(Mux62),
	.datac(temp_imemload_output_201),
	.datad(Mux621),
	.cin(gnd),
	.combout(\temp_rdat_two_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~0 .lut_mask = 16'h4540;
defparam \temp_rdat_two_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N16
cycloneive_lcell_comb \temp_imemload_output~2 (
// Equation(s):
// \temp_imemload_output~2_combout  = (!ex_mem_flush3 & (temp_imemload_output_17 & !use_after_load))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(temp_imemload_output_171),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~2 .lut_mask = 16'h0050;
defparam \temp_imemload_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N18
cycloneive_lcell_comb \temp_imemload_output~3 (
// Equation(s):
// \temp_imemload_output~3_combout  = (temp_imemload_output_16 & (!use_after_load & !ex_mem_flush3))

	.dataa(temp_imemload_output_161),
	.datab(use_after_load),
	.datac(gnd),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_imemload_output~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~3 .lut_mask = 16'h0022;
defparam \temp_imemload_output~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N26
cycloneive_lcell_comb \temp_imemload_output~4 (
// Equation(s):
// \temp_imemload_output~4_combout  = (temp_imemload_output_18 & (!ex_mem_flush3 & !use_after_load))

	.dataa(temp_imemload_output_181),
	.datab(gnd),
	.datac(ex_mem_flush),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~4 .lut_mask = 16'h000A;
defparam \temp_imemload_output~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N16
cycloneive_lcell_comb \temp_imemload_output~5 (
// Equation(s):
// \temp_imemload_output~5_combout  = (temp_imemload_output_19 & (!use_after_load & !ex_mem_flush3))

	.dataa(temp_imemload_output_191),
	.datab(use_after_load),
	.datac(ex_mem_flush),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_imemload_output~5_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~5 .lut_mask = 16'h0202;
defparam \temp_imemload_output~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N16
cycloneive_lcell_comb \temp_imemload_output~6 (
// Equation(s):
// \temp_imemload_output~6_combout  = (!use_after_load & (temp_imemload_output_20 & !ex_mem_flush3))

	.dataa(use_after_load),
	.datab(gnd),
	.datac(temp_imemload_output_201),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_imemload_output~6_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~6 .lut_mask = 16'h0050;
defparam \temp_imemload_output~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N4
cycloneive_lcell_comb \temp_imemload_output~7 (
// Equation(s):
// \temp_imemload_output~7_combout  = (!ex_mem_flush3 & (temp_imemload_output_22 & !use_after_load))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(temp_imemload_output_221),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~7_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~7 .lut_mask = 16'h0030;
defparam \temp_imemload_output~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N26
cycloneive_lcell_comb \temp_imemload_output~8 (
// Equation(s):
// \temp_imemload_output~8_combout  = (temp_imemload_output_21 & (!ex_mem_flush3 & !use_after_load))

	.dataa(temp_imemload_output_211),
	.datab(ex_mem_flush),
	.datac(gnd),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~8_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~8 .lut_mask = 16'h0022;
defparam \temp_imemload_output~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N2
cycloneive_lcell_comb \temp_imemload_output~9 (
// Equation(s):
// \temp_imemload_output~9_combout  = (!use_after_load & (temp_imemload_output_23 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(use_after_load),
	.datac(temp_imemload_output_231),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_imemload_output~9_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~9 .lut_mask = 16'h0030;
defparam \temp_imemload_output~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N4
cycloneive_lcell_comb \temp_imemload_output~10 (
// Equation(s):
// \temp_imemload_output~10_combout  = (!ex_mem_flush3 & (!use_after_load & temp_imemload_output_24))

	.dataa(ex_mem_flush),
	.datab(use_after_load),
	.datac(temp_imemload_output_241),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_imemload_output~10_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~10 .lut_mask = 16'h1010;
defparam \temp_imemload_output~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N16
cycloneive_lcell_comb \temp_imemload_output~11 (
// Equation(s):
// \temp_imemload_output~11_combout  = (!ex_mem_flush3 & (temp_imemload_output_25 & !use_after_load))

	.dataa(ex_mem_flush),
	.datab(temp_imemload_output_251),
	.datac(gnd),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~11_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~11 .lut_mask = 16'h0044;
defparam \temp_imemload_output~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N26
cycloneive_lcell_comb \temp_rdat_one_output~0 (
// Equation(s):
// \temp_rdat_one_output~0_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux301))) # (!temp_imemload_output_25 & (Mux302))))

	.dataa(temp_imemload_output_251),
	.datab(id_ex_flush),
	.datac(Mux301),
	.datad(Mux30),
	.cin(gnd),
	.combout(\temp_rdat_one_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~0 .lut_mask = 16'h3210;
defparam \temp_rdat_one_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N14
cycloneive_lcell_comb \temp_ALUop_output~4 (
// Equation(s):
// \temp_ALUop_output~4_combout  = (extended_imm_16 & ((temp_ALUsrc_output) # ((!temp_imemload_output_31 & WideOr7))))

	.dataa(extended_imm_16),
	.datab(temp_ALUsrc_output),
	.datac(temp_imemload_output_31),
	.datad(WideOr7),
	.cin(gnd),
	.combout(\temp_ALUop_output~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~4 .lut_mask = 16'h8A88;
defparam \temp_ALUop_output~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N20
cycloneive_lcell_comb \temp_ALUop_output~5 (
// Equation(s):
// \temp_ALUop_output~5_combout  = (\temp_ALUsrc_output~0_combout  & temp_imemload_output_5)

	.dataa(gnd),
	.datab(gnd),
	.datac(\temp_ALUsrc_output~0_combout ),
	.datad(temp_imemload_output_51),
	.cin(gnd),
	.combout(\temp_ALUop_output~5_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~5 .lut_mask = 16'hF000;
defparam \temp_ALUop_output~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N16
cycloneive_lcell_comb \temp_ALUop_output~6 (
// Equation(s):
// \temp_ALUop_output~6_combout  = (\temp_ALUop_output~0_combout  & ((\temp_ALUop_output~4_combout ) # ((WideOr1 & \temp_ALUop_output~5_combout ))))

	.dataa(WideOr1),
	.datab(\temp_ALUop_output~0_combout ),
	.datac(\temp_ALUop_output~4_combout ),
	.datad(\temp_ALUop_output~5_combout ),
	.cin(gnd),
	.combout(\temp_ALUop_output~6_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~6 .lut_mask = 16'hC8C0;
defparam \temp_ALUop_output~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N4
cycloneive_lcell_comb \temp_imemload_output~12 (
// Equation(s):
// \temp_imemload_output~12_combout  = (!ex_mem_flush3 & (temp_imemload_output_0 & !use_after_load))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(temp_imemload_output_01),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~12_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~12 .lut_mask = 16'h0050;
defparam \temp_imemload_output~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N26
cycloneive_lcell_comb \temp_imemload_output~13 (
// Equation(s):
// \temp_imemload_output~13_combout  = (!ex_mem_flush3 & (!use_after_load & temp_imemload_output_6))

	.dataa(ex_mem_flush),
	.datab(use_after_load),
	.datac(gnd),
	.datad(temp_imemload_output_61),
	.cin(gnd),
	.combout(\temp_imemload_output~13_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~13 .lut_mask = 16'h1100;
defparam \temp_imemload_output~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N4
cycloneive_lcell_comb \temp_rdat_two_output~1 (
// Equation(s):
// \temp_rdat_two_output~1_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux63)) # (!temp_imemload_output_20 & ((Mux631)))))

	.dataa(Mux63),
	.datab(id_ex_flush),
	.datac(temp_imemload_output_201),
	.datad(Mux631),
	.cin(gnd),
	.combout(\temp_rdat_two_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~1 .lut_mask = 16'h2320;
defparam \temp_rdat_two_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N28
cycloneive_lcell_comb \temp_rdat_one_output~1 (
// Equation(s):
// \temp_rdat_one_output~1_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux311))) # (!temp_imemload_output_25 & (Mux312))))

	.dataa(temp_imemload_output_251),
	.datab(id_ex_flush),
	.datac(Mux311),
	.datad(Mux31),
	.cin(gnd),
	.combout(\temp_rdat_one_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~1 .lut_mask = 16'h3210;
defparam \temp_rdat_one_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N30
cycloneive_lcell_comb \temp_rdat_one_output~2 (
// Equation(s):
// \temp_rdat_one_output~2_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux291)) # (!temp_imemload_output_25 & ((Mux292)))))

	.dataa(Mux29),
	.datab(id_ex_flush),
	.datac(Mux291),
	.datad(temp_imemload_output_251),
	.cin(gnd),
	.combout(\temp_rdat_one_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~2 .lut_mask = 16'h2230;
defparam \temp_rdat_one_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N0
cycloneive_lcell_comb \temp_rdat_one_output~3 (
// Equation(s):
// \temp_rdat_one_output~3_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux271)) # (!temp_imemload_output_25 & ((Mux272)))))

	.dataa(Mux27),
	.datab(id_ex_flush),
	.datac(temp_imemload_output_251),
	.datad(Mux271),
	.cin(gnd),
	.combout(\temp_rdat_one_output~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~3 .lut_mask = 16'h2320;
defparam \temp_rdat_one_output~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N18
cycloneive_lcell_comb \temp_rdat_one_output~4 (
// Equation(s):
// \temp_rdat_one_output~4_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux281))) # (!temp_imemload_output_25 & (Mux282))))

	.dataa(Mux281),
	.datab(temp_imemload_output_251),
	.datac(id_ex_flush),
	.datad(Mux28),
	.cin(gnd),
	.combout(\temp_rdat_one_output~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~4 .lut_mask = 16'h0E02;
defparam \temp_rdat_one_output~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N28
cycloneive_lcell_comb \temp_imemload_output~14 (
// Equation(s):
// \temp_imemload_output~14_combout  = (!ex_mem_flush3 & (!use_after_load & temp_imemload_output_2))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(use_after_load),
	.datad(temp_imemload_output_210),
	.cin(gnd),
	.combout(\temp_imemload_output~14_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~14 .lut_mask = 16'h0300;
defparam \temp_imemload_output~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N16
cycloneive_lcell_comb \temp_imemload_output~15 (
// Equation(s):
// \temp_imemload_output~15_combout  = (!ex_mem_flush3 & (!use_after_load & temp_imemload_output_8))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(use_after_load),
	.datad(temp_imemload_output_81),
	.cin(gnd),
	.combout(\temp_imemload_output~15_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~15 .lut_mask = 16'h0500;
defparam \temp_imemload_output~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N28
cycloneive_lcell_comb \temp_rdat_two_output~2 (
// Equation(s):
// \temp_rdat_two_output~2_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux61))) # (!temp_imemload_output_20 & (Mux611))))

	.dataa(Mux611),
	.datab(Mux61),
	.datac(id_ex_flush),
	.datad(temp_imemload_output_201),
	.cin(gnd),
	.combout(\temp_rdat_two_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~2 .lut_mask = 16'h0C0A;
defparam \temp_rdat_two_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N8
cycloneive_lcell_comb \temp_rdat_one_output~5 (
// Equation(s):
// \temp_rdat_one_output~5_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux231)) # (!temp_imemload_output_25 & ((Mux232)))))

	.dataa(Mux23),
	.datab(id_ex_flush),
	.datac(temp_imemload_output_251),
	.datad(Mux231),
	.cin(gnd),
	.combout(\temp_rdat_one_output~5_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~5 .lut_mask = 16'h2320;
defparam \temp_rdat_one_output~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N24
cycloneive_lcell_comb \temp_rdat_one_output~6 (
// Equation(s):
// \temp_rdat_one_output~6_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux241)) # (!temp_imemload_output_25 & ((Mux242)))))

	.dataa(Mux24),
	.datab(id_ex_flush),
	.datac(temp_imemload_output_251),
	.datad(Mux241),
	.cin(gnd),
	.combout(\temp_rdat_one_output~6_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~6 .lut_mask = 16'h2320;
defparam \temp_rdat_one_output~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N26
cycloneive_lcell_comb \temp_rdat_one_output~7 (
// Equation(s):
// \temp_rdat_one_output~7_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux251)) # (!temp_imemload_output_25 & ((Mux252)))))

	.dataa(Mux25),
	.datab(temp_imemload_output_251),
	.datac(id_ex_flush),
	.datad(Mux251),
	.cin(gnd),
	.combout(\temp_rdat_one_output~7_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~7 .lut_mask = 16'h0B08;
defparam \temp_rdat_one_output~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N14
cycloneive_lcell_comb \temp_rdat_one_output~8 (
// Equation(s):
// \temp_rdat_one_output~8_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux261))) # (!temp_imemload_output_25 & (Mux262))))

	.dataa(temp_imemload_output_251),
	.datab(id_ex_flush),
	.datac(Mux261),
	.datad(Mux26),
	.cin(gnd),
	.combout(\temp_rdat_one_output~8_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~8 .lut_mask = 16'h3210;
defparam \temp_rdat_one_output~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N26
cycloneive_lcell_comb \temp_imemload_output~16 (
// Equation(s):
// \temp_imemload_output~16_combout  = (!ex_mem_flush3 & (!use_after_load & temp_imemload_output_3))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(use_after_load),
	.datad(temp_imemload_output_32),
	.cin(gnd),
	.combout(\temp_imemload_output~16_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~16 .lut_mask = 16'h0500;
defparam \temp_imemload_output~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N8
cycloneive_lcell_comb \temp_imemload_output~17 (
// Equation(s):
// \temp_imemload_output~17_combout  = (!ex_mem_flush3 & (!use_after_load & temp_imemload_output_9))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(use_after_load),
	.datad(temp_imemload_output_91),
	.cin(gnd),
	.combout(\temp_imemload_output~17_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~17 .lut_mask = 16'h0500;
defparam \temp_imemload_output~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N16
cycloneive_lcell_comb \temp_rdat_two_output~3 (
// Equation(s):
// \temp_rdat_two_output~3_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux60))) # (!temp_imemload_output_20 & (Mux601))))

	.dataa(id_ex_flush),
	.datab(temp_imemload_output_201),
	.datac(Mux601),
	.datad(Mux60),
	.cin(gnd),
	.combout(\temp_rdat_two_output~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~3 .lut_mask = 16'h5410;
defparam \temp_rdat_two_output~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N0
cycloneive_lcell_comb \temp_rdat_one_output~9 (
// Equation(s):
// \temp_rdat_one_output~9_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux151))) # (!temp_imemload_output_25 & (Mux152))))

	.dataa(Mux151),
	.datab(Mux15),
	.datac(temp_imemload_output_251),
	.datad(id_ex_flush),
	.cin(gnd),
	.combout(\temp_rdat_one_output~9_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~9 .lut_mask = 16'h00CA;
defparam \temp_rdat_one_output~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N24
cycloneive_lcell_comb \temp_rdat_one_output~10 (
// Equation(s):
// \temp_rdat_one_output~10_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux171))) # (!temp_imemload_output_25 & (Mux172))))

	.dataa(Mux171),
	.datab(temp_imemload_output_251),
	.datac(Mux17),
	.datad(id_ex_flush),
	.cin(gnd),
	.combout(\temp_rdat_one_output~10_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~10 .lut_mask = 16'h00E2;
defparam \temp_rdat_one_output~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N22
cycloneive_lcell_comb \temp_rdat_one_output~11 (
// Equation(s):
// \temp_rdat_one_output~11_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux161)) # (!temp_imemload_output_25 & ((Mux162)))))

	.dataa(id_ex_flush),
	.datab(Mux16),
	.datac(Mux161),
	.datad(temp_imemload_output_251),
	.cin(gnd),
	.combout(\temp_rdat_one_output~11_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~11 .lut_mask = 16'h4450;
defparam \temp_rdat_one_output~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N30
cycloneive_lcell_comb \temp_rdat_one_output~12 (
// Equation(s):
// \temp_rdat_one_output~12_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux181)) # (!temp_imemload_output_25 & ((Mux182)))))

	.dataa(Mux18),
	.datab(id_ex_flush),
	.datac(temp_imemload_output_251),
	.datad(Mux181),
	.cin(gnd),
	.combout(\temp_rdat_one_output~12_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~12 .lut_mask = 16'h2320;
defparam \temp_rdat_one_output~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y43_N24
cycloneive_lcell_comb \temp_rdat_one_output~13 (
// Equation(s):
// \temp_rdat_one_output~13_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux191))) # (!temp_imemload_output_25 & (Mux192))))

	.dataa(id_ex_flush),
	.datab(Mux191),
	.datac(temp_imemload_output_251),
	.datad(Mux19),
	.cin(gnd),
	.combout(\temp_rdat_one_output~13_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~13 .lut_mask = 16'h5404;
defparam \temp_rdat_one_output~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N30
cycloneive_lcell_comb \temp_rdat_one_output~14 (
// Equation(s):
// \temp_rdat_one_output~14_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux211)) # (!temp_imemload_output_25 & ((Mux212)))))

	.dataa(temp_imemload_output_251),
	.datab(id_ex_flush),
	.datac(Mux21),
	.datad(Mux211),
	.cin(gnd),
	.combout(\temp_rdat_one_output~14_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~14 .lut_mask = 16'h3120;
defparam \temp_rdat_one_output~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N14
cycloneive_lcell_comb \temp_rdat_one_output~15 (
// Equation(s):
// \temp_rdat_one_output~15_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux201)) # (!temp_imemload_output_25 & ((Mux202)))))

	.dataa(temp_imemload_output_251),
	.datab(Mux20),
	.datac(Mux201),
	.datad(id_ex_flush),
	.cin(gnd),
	.combout(\temp_rdat_one_output~15_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~15 .lut_mask = 16'h00D8;
defparam \temp_rdat_one_output~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N18
cycloneive_lcell_comb \temp_rdat_one_output~16 (
// Equation(s):
// \temp_rdat_one_output~16_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux221))) # (!temp_imemload_output_25 & (Mux222))))

	.dataa(Mux221),
	.datab(Mux22),
	.datac(id_ex_flush),
	.datad(temp_imemload_output_251),
	.cin(gnd),
	.combout(\temp_rdat_one_output~16_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~16 .lut_mask = 16'h0C0A;
defparam \temp_rdat_one_output~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N28
cycloneive_lcell_comb \temp_imemload_output~18 (
// Equation(s):
// \temp_imemload_output~18_combout  = (!ex_mem_flush3 & (temp_imemload_output_4 & !use_after_load))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(temp_imemload_output_41),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~18_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~18 .lut_mask = 16'h0050;
defparam \temp_imemload_output~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N22
cycloneive_lcell_comb \temp_imemload_output~19 (
// Equation(s):
// \temp_imemload_output~19_combout  = (!use_after_load & (!ex_mem_flush3 & temp_imemload_output_10))

	.dataa(use_after_load),
	.datab(ex_mem_flush),
	.datac(gnd),
	.datad(temp_imemload_output_101),
	.cin(gnd),
	.combout(\temp_imemload_output~19_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~19 .lut_mask = 16'h1100;
defparam \temp_imemload_output~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N16
cycloneive_lcell_comb \temp_rdat_two_output~4 (
// Equation(s):
// \temp_rdat_two_output~4_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux59)) # (!temp_imemload_output_20 & ((Mux591)))))

	.dataa(Mux59),
	.datab(id_ex_flush),
	.datac(temp_imemload_output_201),
	.datad(Mux591),
	.cin(gnd),
	.combout(\temp_rdat_two_output~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~4 .lut_mask = 16'h2320;
defparam \temp_rdat_two_output~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N2
cycloneive_lcell_comb \temp_rdat_one_output~17 (
// Equation(s):
// \temp_rdat_one_output~17_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux01)) # (!temp_imemload_output_25 & ((Mux02)))))

	.dataa(temp_imemload_output_251),
	.datab(Mux0),
	.datac(id_ex_flush),
	.datad(Mux01),
	.cin(gnd),
	.combout(\temp_rdat_one_output~17_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~17 .lut_mask = 16'h0D08;
defparam \temp_rdat_one_output~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N2
cycloneive_lcell_comb \temp_rdat_one_output~18 (
// Equation(s):
// \temp_rdat_one_output~18_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux110)) # (!temp_imemload_output_25 & ((Mux111)))))

	.dataa(id_ex_flush),
	.datab(Mux1),
	.datac(Mux11),
	.datad(temp_imemload_output_251),
	.cin(gnd),
	.combout(\temp_rdat_one_output~18_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~18 .lut_mask = 16'h4450;
defparam \temp_rdat_one_output~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N0
cycloneive_lcell_comb \temp_rdat_one_output~19 (
// Equation(s):
// \temp_rdat_one_output~19_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux210)) # (!temp_imemload_output_25 & ((Mux213)))))

	.dataa(Mux2),
	.datab(id_ex_flush),
	.datac(Mux210),
	.datad(temp_imemload_output_251),
	.cin(gnd),
	.combout(\temp_rdat_one_output~19_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~19 .lut_mask = 16'h2230;
defparam \temp_rdat_one_output~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N28
cycloneive_lcell_comb \temp_rdat_one_output~20 (
// Equation(s):
// \temp_rdat_one_output~20_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux51)) # (!temp_imemload_output_25 & ((Mux52)))))

	.dataa(id_ex_flush),
	.datab(Mux5),
	.datac(temp_imemload_output_251),
	.datad(Mux51),
	.cin(gnd),
	.combout(\temp_rdat_one_output~20_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~20 .lut_mask = 16'h4540;
defparam \temp_rdat_one_output~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N0
cycloneive_lcell_comb \temp_rdat_one_output~21 (
// Equation(s):
// \temp_rdat_one_output~21_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux64))) # (!temp_imemload_output_25 & (Mux65))))

	.dataa(id_ex_flush),
	.datab(Mux64),
	.datac(temp_imemload_output_251),
	.datad(Mux6),
	.cin(gnd),
	.combout(\temp_rdat_one_output~21_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~21 .lut_mask = 16'h5404;
defparam \temp_rdat_one_output~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N12
cycloneive_lcell_comb \temp_rdat_one_output~22 (
// Equation(s):
// \temp_rdat_one_output~22_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux32))) # (!temp_imemload_output_25 & (Mux33))))

	.dataa(id_ex_flush),
	.datab(temp_imemload_output_251),
	.datac(Mux32),
	.datad(Mux3),
	.cin(gnd),
	.combout(\temp_rdat_one_output~22_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~22 .lut_mask = 16'h5410;
defparam \temp_rdat_one_output~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N0
cycloneive_lcell_comb \temp_rdat_one_output~23 (
// Equation(s):
// \temp_rdat_one_output~23_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux41)) # (!temp_imemload_output_25 & ((Mux42)))))

	.dataa(id_ex_flush),
	.datab(Mux4),
	.datac(Mux41),
	.datad(temp_imemload_output_251),
	.cin(gnd),
	.combout(\temp_rdat_one_output~23_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~23 .lut_mask = 16'h4450;
defparam \temp_rdat_one_output~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N8
cycloneive_lcell_comb \temp_rdat_one_output~24 (
// Equation(s):
// \temp_rdat_one_output~24_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux141)) # (!temp_imemload_output_25 & ((Mux142)))))

	.dataa(Mux14),
	.datab(Mux141),
	.datac(temp_imemload_output_251),
	.datad(id_ex_flush),
	.cin(gnd),
	.combout(\temp_rdat_one_output~24_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~24 .lut_mask = 16'h00AC;
defparam \temp_rdat_one_output~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N10
cycloneive_lcell_comb \temp_rdat_one_output~25 (
// Equation(s):
// \temp_rdat_one_output~25_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux112))) # (!temp_imemload_output_25 & (Mux113))))

	.dataa(id_ex_flush),
	.datab(Mux112),
	.datac(temp_imemload_output_251),
	.datad(Mux111),
	.cin(gnd),
	.combout(\temp_rdat_one_output~25_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~25 .lut_mask = 16'h5404;
defparam \temp_rdat_one_output~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N10
cycloneive_lcell_comb \temp_rdat_one_output~26 (
// Equation(s):
// \temp_rdat_one_output~26_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux121)) # (!temp_imemload_output_25 & ((Mux122)))))

	.dataa(temp_imemload_output_251),
	.datab(id_ex_flush),
	.datac(Mux12),
	.datad(Mux121),
	.cin(gnd),
	.combout(\temp_rdat_one_output~26_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~26 .lut_mask = 16'h3120;
defparam \temp_rdat_one_output~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N14
cycloneive_lcell_comb \temp_rdat_one_output~27 (
// Equation(s):
// \temp_rdat_one_output~27_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux131))) # (!temp_imemload_output_25 & (Mux132))))

	.dataa(id_ex_flush),
	.datab(Mux131),
	.datac(Mux13),
	.datad(temp_imemload_output_251),
	.cin(gnd),
	.combout(\temp_rdat_one_output~27_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~27 .lut_mask = 16'h5044;
defparam \temp_rdat_one_output~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N14
cycloneive_lcell_comb \temp_rdat_one_output~28 (
// Equation(s):
// \temp_rdat_one_output~28_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux71))) # (!temp_imemload_output_25 & (Mux72))))

	.dataa(temp_imemload_output_251),
	.datab(Mux71),
	.datac(Mux7),
	.datad(id_ex_flush),
	.cin(gnd),
	.combout(\temp_rdat_one_output~28_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~28 .lut_mask = 16'h00E4;
defparam \temp_rdat_one_output~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N16
cycloneive_lcell_comb \temp_rdat_one_output~29 (
// Equation(s):
// \temp_rdat_one_output~29_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux81))) # (!temp_imemload_output_25 & (Mux82))))

	.dataa(Mux81),
	.datab(temp_imemload_output_251),
	.datac(Mux8),
	.datad(id_ex_flush),
	.cin(gnd),
	.combout(\temp_rdat_one_output~29_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~29 .lut_mask = 16'h00E2;
defparam \temp_rdat_one_output~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N24
cycloneive_lcell_comb \temp_rdat_one_output~30 (
// Equation(s):
// \temp_rdat_one_output~30_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & (Mux91)) # (!temp_imemload_output_25 & ((Mux92)))))

	.dataa(Mux9),
	.datab(Mux91),
	.datac(temp_imemload_output_251),
	.datad(id_ex_flush),
	.cin(gnd),
	.combout(\temp_rdat_one_output~30_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~30 .lut_mask = 16'h00AC;
defparam \temp_rdat_one_output~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N14
cycloneive_lcell_comb \temp_rdat_one_output~31 (
// Equation(s):
// \temp_rdat_one_output~31_combout  = (!id_ex_flush1 & ((temp_imemload_output_25 & ((Mux101))) # (!temp_imemload_output_25 & (Mux102))))

	.dataa(Mux101),
	.datab(temp_imemload_output_251),
	.datac(id_ex_flush),
	.datad(Mux10),
	.cin(gnd),
	.combout(\temp_rdat_one_output~31_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_one_output~31 .lut_mask = 16'h0E02;
defparam \temp_rdat_one_output~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N18
cycloneive_lcell_comb \temp_rdat_two_output~5 (
// Equation(s):
// \temp_rdat_two_output~5_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux48)) # (!temp_imemload_output_20 & ((Mux481)))))

	.dataa(Mux48),
	.datab(temp_imemload_output_201),
	.datac(Mux481),
	.datad(id_ex_flush),
	.cin(gnd),
	.combout(\temp_rdat_two_output~5_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~5 .lut_mask = 16'h00B8;
defparam \temp_rdat_two_output~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N6
cycloneive_lcell_comb \temp_imemload_output~20 (
// Equation(s):
// \temp_imemload_output~20_combout  = (!use_after_load & (!ex_mem_flush3 & temp_imemload_output_15))

	.dataa(gnd),
	.datab(use_after_load),
	.datac(ex_mem_flush),
	.datad(temp_imemload_output_151),
	.cin(gnd),
	.combout(\temp_imemload_output~20_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~20 .lut_mask = 16'h0300;
defparam \temp_imemload_output~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N4
cycloneive_lcell_comb \temp_rdat_two_output~6 (
// Equation(s):
// \temp_rdat_two_output~6_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux511))) # (!temp_imemload_output_20 & (Mux512))))

	.dataa(temp_imemload_output_201),
	.datab(Mux512),
	.datac(id_ex_flush),
	.datad(Mux511),
	.cin(gnd),
	.combout(\temp_rdat_two_output~6_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~6 .lut_mask = 16'h0E04;
defparam \temp_rdat_two_output~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N26
cycloneive_lcell_comb \temp_imemload_output~21 (
// Equation(s):
// \temp_imemload_output~21_combout  = (!ex_mem_flush3 & (!use_after_load & temp_imemload_output_12))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(use_after_load),
	.datad(temp_imemload_output_121),
	.cin(gnd),
	.combout(\temp_imemload_output~21_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~21 .lut_mask = 16'h0300;
defparam \temp_imemload_output~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N12
cycloneive_lcell_comb \temp_rdat_two_output~7 (
// Equation(s):
// \temp_rdat_two_output~7_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux36))) # (!temp_imemload_output_20 & (Mux361))))

	.dataa(id_ex_flush),
	.datab(Mux361),
	.datac(temp_imemload_output_201),
	.datad(Mux36),
	.cin(gnd),
	.combout(\temp_rdat_two_output~7_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~7 .lut_mask = 16'h5404;
defparam \temp_rdat_two_output~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N4
cycloneive_lcell_comb \temp_rdat_two_output~8 (
// Equation(s):
// \temp_rdat_two_output~8_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux45)) # (!temp_imemload_output_20 & ((Mux451)))))

	.dataa(id_ex_flush),
	.datab(Mux45),
	.datac(Mux451),
	.datad(temp_imemload_output_201),
	.cin(gnd),
	.combout(\temp_rdat_two_output~8_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~8 .lut_mask = 16'h4450;
defparam \temp_rdat_two_output~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N22
cycloneive_lcell_comb \temp_rdat_two_output~9 (
// Equation(s):
// \temp_rdat_two_output~9_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux46))) # (!temp_imemload_output_20 & (Mux461))))

	.dataa(Mux461),
	.datab(Mux46),
	.datac(temp_imemload_output_201),
	.datad(id_ex_flush),
	.cin(gnd),
	.combout(\temp_rdat_two_output~9_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~9 .lut_mask = 16'h00CA;
defparam \temp_rdat_two_output~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N2
cycloneive_lcell_comb \temp_rdat_two_output~10 (
// Equation(s):
// \temp_rdat_two_output~10_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux47))) # (!temp_imemload_output_20 & (Mux471))))

	.dataa(temp_imemload_output_201),
	.datab(id_ex_flush),
	.datac(Mux471),
	.datad(Mux47),
	.cin(gnd),
	.combout(\temp_rdat_two_output~10_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~10 .lut_mask = 16'h3210;
defparam \temp_rdat_two_output~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N22
cycloneive_lcell_comb \temp_rdat_two_output~11 (
// Equation(s):
// \temp_rdat_two_output~11_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux321)) # (!temp_imemload_output_20 & ((Mux322)))))

	.dataa(Mux321),
	.datab(Mux322),
	.datac(id_ex_flush),
	.datad(temp_imemload_output_201),
	.cin(gnd),
	.combout(\temp_rdat_two_output~11_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~11 .lut_mask = 16'h0A0C;
defparam \temp_rdat_two_output~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N30
cycloneive_lcell_comb \temp_rdat_two_output~12 (
// Equation(s):
// \temp_rdat_two_output~12_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux331)) # (!temp_imemload_output_20 & ((Mux332)))))

	.dataa(id_ex_flush),
	.datab(Mux33),
	.datac(Mux331),
	.datad(temp_imemload_output_201),
	.cin(gnd),
	.combout(\temp_rdat_two_output~12_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~12 .lut_mask = 16'h4450;
defparam \temp_rdat_two_output~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N12
cycloneive_lcell_comb \temp_rdat_two_output~13 (
// Equation(s):
// \temp_rdat_two_output~13_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux34))) # (!temp_imemload_output_20 & (Mux341))))

	.dataa(temp_imemload_output_201),
	.datab(Mux341),
	.datac(id_ex_flush),
	.datad(Mux34),
	.cin(gnd),
	.combout(\temp_rdat_two_output~13_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~13 .lut_mask = 16'h0E04;
defparam \temp_rdat_two_output~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N4
cycloneive_lcell_comb \temp_rdat_two_output~14 (
// Equation(s):
// \temp_rdat_two_output~14_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux35))) # (!temp_imemload_output_20 & (Mux351))))

	.dataa(temp_imemload_output_201),
	.datab(Mux351),
	.datac(id_ex_flush),
	.datad(Mux35),
	.cin(gnd),
	.combout(\temp_rdat_two_output~14_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~14 .lut_mask = 16'h0E04;
defparam \temp_rdat_two_output~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N24
cycloneive_lcell_comb \temp_rdat_two_output~15 (
// Equation(s):
// \temp_rdat_two_output~15_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux37)) # (!temp_imemload_output_20 & ((Mux371)))))

	.dataa(id_ex_flush),
	.datab(temp_imemload_output_201),
	.datac(Mux37),
	.datad(Mux371),
	.cin(gnd),
	.combout(\temp_rdat_two_output~15_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~15 .lut_mask = 16'h5140;
defparam \temp_rdat_two_output~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N14
cycloneive_lcell_comb \temp_rdat_two_output~16 (
// Equation(s):
// \temp_rdat_two_output~16_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux38)) # (!temp_imemload_output_20 & ((Mux381)))))

	.dataa(temp_imemload_output_201),
	.datab(id_ex_flush),
	.datac(Mux38),
	.datad(Mux381),
	.cin(gnd),
	.combout(\temp_rdat_two_output~16_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~16 .lut_mask = 16'h3120;
defparam \temp_rdat_two_output~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N28
cycloneive_lcell_comb \temp_rdat_two_output~17 (
// Equation(s):
// \temp_rdat_two_output~17_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux39)) # (!temp_imemload_output_20 & ((Mux391)))))

	.dataa(Mux39),
	.datab(Mux391),
	.datac(temp_imemload_output_201),
	.datad(id_ex_flush),
	.cin(gnd),
	.combout(\temp_rdat_two_output~17_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~17 .lut_mask = 16'h00AC;
defparam \temp_rdat_two_output~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N4
cycloneive_lcell_comb \temp_rdat_two_output~18 (
// Equation(s):
// \temp_rdat_two_output~18_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux40)) # (!temp_imemload_output_20 & ((Mux401)))))

	.dataa(temp_imemload_output_201),
	.datab(Mux40),
	.datac(id_ex_flush),
	.datad(Mux401),
	.cin(gnd),
	.combout(\temp_rdat_two_output~18_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~18 .lut_mask = 16'h0D08;
defparam \temp_rdat_two_output~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N2
cycloneive_lcell_comb \temp_rdat_two_output~19 (
// Equation(s):
// \temp_rdat_two_output~19_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux411))) # (!temp_imemload_output_20 & (Mux412))))

	.dataa(temp_imemload_output_201),
	.datab(Mux412),
	.datac(id_ex_flush),
	.datad(Mux411),
	.cin(gnd),
	.combout(\temp_rdat_two_output~19_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~19 .lut_mask = 16'h0E04;
defparam \temp_rdat_two_output~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N24
cycloneive_lcell_comb \temp_rdat_two_output~20 (
// Equation(s):
// \temp_rdat_two_output~20_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux421))) # (!temp_imemload_output_20 & (Mux422))))

	.dataa(Mux421),
	.datab(temp_imemload_output_201),
	.datac(id_ex_flush),
	.datad(Mux42),
	.cin(gnd),
	.combout(\temp_rdat_two_output~20_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~20 .lut_mask = 16'h0E02;
defparam \temp_rdat_two_output~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N16
cycloneive_lcell_comb \temp_rdat_two_output~21 (
// Equation(s):
// \temp_rdat_two_output~21_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux43)) # (!temp_imemload_output_20 & ((Mux431)))))

	.dataa(id_ex_flush),
	.datab(Mux43),
	.datac(temp_imemload_output_201),
	.datad(Mux431),
	.cin(gnd),
	.combout(\temp_rdat_two_output~21_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~21 .lut_mask = 16'h4540;
defparam \temp_rdat_two_output~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N28
cycloneive_lcell_comb \temp_rdat_two_output~22 (
// Equation(s):
// \temp_rdat_two_output~22_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux44))) # (!temp_imemload_output_20 & (Mux441))))

	.dataa(id_ex_flush),
	.datab(temp_imemload_output_201),
	.datac(Mux441),
	.datad(Mux44),
	.cin(gnd),
	.combout(\temp_rdat_two_output~22_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~22 .lut_mask = 16'h5410;
defparam \temp_rdat_two_output~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N20
cycloneive_lcell_comb \temp_imemload_output~22 (
// Equation(s):
// \temp_imemload_output~22_combout  = (temp_imemload_output_14 & (!use_after_load & !ex_mem_flush3))

	.dataa(temp_imemload_output_141),
	.datab(use_after_load),
	.datac(ex_mem_flush),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_imemload_output~22_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~22 .lut_mask = 16'h0202;
defparam \temp_imemload_output~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N20
cycloneive_lcell_comb \temp_rdat_two_output~23 (
// Equation(s):
// \temp_rdat_two_output~23_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux53)) # (!temp_imemload_output_20 & ((Mux531)))))

	.dataa(Mux53),
	.datab(id_ex_flush),
	.datac(Mux531),
	.datad(temp_imemload_output_201),
	.cin(gnd),
	.combout(\temp_rdat_two_output~23_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~23 .lut_mask = 16'h2230;
defparam \temp_rdat_two_output~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N12
cycloneive_lcell_comb \temp_rdat_two_output~24 (
// Equation(s):
// \temp_rdat_two_output~24_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux49))) # (!temp_imemload_output_20 & (Mux491))))

	.dataa(id_ex_flush),
	.datab(Mux491),
	.datac(temp_imemload_output_201),
	.datad(Mux49),
	.cin(gnd),
	.combout(\temp_rdat_two_output~24_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~24 .lut_mask = 16'h5404;
defparam \temp_rdat_two_output~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N12
cycloneive_lcell_comb \temp_rdat_two_output~25 (
// Equation(s):
// \temp_rdat_two_output~25_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux54)) # (!temp_imemload_output_20 & ((Mux541)))))

	.dataa(temp_imemload_output_201),
	.datab(id_ex_flush),
	.datac(Mux54),
	.datad(Mux541),
	.cin(gnd),
	.combout(\temp_rdat_two_output~25_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~25 .lut_mask = 16'h3120;
defparam \temp_rdat_two_output~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N6
cycloneive_lcell_comb \temp_rdat_two_output~26 (
// Equation(s):
// \temp_rdat_two_output~26_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux55))) # (!temp_imemload_output_20 & (Mux551))))

	.dataa(temp_imemload_output_201),
	.datab(Mux551),
	.datac(id_ex_flush),
	.datad(Mux55),
	.cin(gnd),
	.combout(\temp_rdat_two_output~26_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~26 .lut_mask = 16'h0E04;
defparam \temp_rdat_two_output~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N18
cycloneive_lcell_comb \temp_rdat_two_output~27 (
// Equation(s):
// \temp_rdat_two_output~27_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux56)) # (!temp_imemload_output_20 & ((Mux561)))))

	.dataa(Mux56),
	.datab(id_ex_flush),
	.datac(Mux561),
	.datad(temp_imemload_output_201),
	.cin(gnd),
	.combout(\temp_rdat_two_output~27_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~27 .lut_mask = 16'h2230;
defparam \temp_rdat_two_output~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N16
cycloneive_lcell_comb \temp_rdat_two_output~28 (
// Equation(s):
// \temp_rdat_two_output~28_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux57))) # (!temp_imemload_output_20 & (Mux571))))

	.dataa(temp_imemload_output_201),
	.datab(Mux571),
	.datac(id_ex_flush),
	.datad(Mux57),
	.cin(gnd),
	.combout(\temp_rdat_two_output~28_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~28 .lut_mask = 16'h0E04;
defparam \temp_rdat_two_output~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N20
cycloneive_lcell_comb \temp_rdat_two_output~29 (
// Equation(s):
// \temp_rdat_two_output~29_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux58))) # (!temp_imemload_output_20 & (Mux581))))

	.dataa(temp_imemload_output_201),
	.datab(id_ex_flush),
	.datac(Mux581),
	.datad(Mux58),
	.cin(gnd),
	.combout(\temp_rdat_two_output~29_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~29 .lut_mask = 16'h3210;
defparam \temp_rdat_two_output~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N30
cycloneive_lcell_comb \temp_imemload_output~23 (
// Equation(s):
// \temp_imemload_output~23_combout  = (temp_imemload_output_5 & (!use_after_load & !ex_mem_flush3))

	.dataa(temp_imemload_output_51),
	.datab(use_after_load),
	.datac(gnd),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_imemload_output~23_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~23 .lut_mask = 16'h0022;
defparam \temp_imemload_output~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N10
cycloneive_lcell_comb \temp_rdat_two_output~30 (
// Equation(s):
// \temp_rdat_two_output~30_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & ((Mux50))) # (!temp_imemload_output_20 & (Mux501))))

	.dataa(Mux501),
	.datab(id_ex_flush),
	.datac(temp_imemload_output_201),
	.datad(Mux50),
	.cin(gnd),
	.combout(\temp_rdat_two_output~30_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~30 .lut_mask = 16'h3202;
defparam \temp_rdat_two_output~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N20
cycloneive_lcell_comb \temp_imemload_output~24 (
// Equation(s):
// \temp_imemload_output~24_combout  = (!ex_mem_flush3 & (!use_after_load & temp_imemload_output_13))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(use_after_load),
	.datad(temp_imemload_output_131),
	.cin(gnd),
	.combout(\temp_imemload_output~24_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~24 .lut_mask = 16'h0500;
defparam \temp_imemload_output~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N30
cycloneive_lcell_comb \temp_rdat_two_output~31 (
// Equation(s):
// \temp_rdat_two_output~31_combout  = (!id_ex_flush1 & ((temp_imemload_output_20 & (Mux521)) # (!temp_imemload_output_20 & ((Mux522)))))

	.dataa(id_ex_flush),
	.datab(Mux52),
	.datac(Mux521),
	.datad(temp_imemload_output_201),
	.cin(gnd),
	.combout(\temp_rdat_two_output~31_combout ),
	.cout());
// synopsys translate_off
defparam \temp_rdat_two_output~31 .lut_mask = 16'h4450;
defparam \temp_rdat_two_output~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N24
cycloneive_lcell_comb \temp_imemload_output~25 (
// Equation(s):
// \temp_imemload_output~25_combout  = (!ex_mem_flush3 & (!use_after_load & temp_imemload_output_11))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(use_after_load),
	.datad(temp_imemload_output_111),
	.cin(gnd),
	.combout(\temp_imemload_output~25_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~25 .lut_mask = 16'h0300;
defparam \temp_imemload_output~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N18
cycloneive_lcell_comb \temp_ALUop_output~7 (
// Equation(s):
// \temp_ALUop_output~7_combout  = (extended_imm_16 & ((temp_ALUsrc_output) # ((WideOr6 & !temp_imemload_output_31))))

	.dataa(extended_imm_16),
	.datab(WideOr6),
	.datac(temp_imemload_output_31),
	.datad(temp_ALUsrc_output),
	.cin(gnd),
	.combout(\temp_ALUop_output~7_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~7 .lut_mask = 16'hAA08;
defparam \temp_ALUop_output~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N10
cycloneive_lcell_comb \temp_ALUop_output~8 (
// Equation(s):
// \temp_ALUop_output~8_combout  = (\temp_ALUop_output~0_combout  & ((\temp_ALUop_output~7_combout ) # ((WideOr0 & \temp_ALUop_output~5_combout ))))

	.dataa(WideOr0),
	.datab(\temp_ALUop_output~5_combout ),
	.datac(\temp_ALUop_output~0_combout ),
	.datad(\temp_ALUop_output~7_combout ),
	.cin(gnd),
	.combout(\temp_ALUop_output~8_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~8 .lut_mask = 16'hF080;
defparam \temp_ALUop_output~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N2
cycloneive_lcell_comb \temp_ALUop_output~9 (
// Equation(s):
// \temp_ALUop_output~9_combout  = (halt_out & (!temp_imemload_output_2 & \temp_ALUsrc_output~0_combout ))

	.dataa(halt_out),
	.datab(temp_imemload_output_210),
	.datac(\temp_ALUsrc_output~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_ALUop_output~9_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~9 .lut_mask = 16'h2020;
defparam \temp_ALUop_output~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N16
cycloneive_lcell_comb \temp_ALUop_output~10 (
// Equation(s):
// \temp_ALUop_output~10_combout  = (!temp_imemload_output_30 & (!temp_imemload_output_31 & (temp_imemload_output_29 & !temp_imemload_output_28)))

	.dataa(temp_imemload_output_30),
	.datab(temp_imemload_output_31),
	.datac(temp_imemload_output_29),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(\temp_ALUop_output~10_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~10 .lut_mask = 16'h0010;
defparam \temp_ALUop_output~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N28
cycloneive_lcell_comb \temp_ALUop_output~11 (
// Equation(s):
// \temp_ALUop_output~11_combout  = (\temp_ALUop_output~0_combout  & ((\temp_ALUop_output~9_combout ) # ((temp_imemload_output_27 & \temp_ALUop_output~10_combout ))))

	.dataa(\temp_ALUop_output~9_combout ),
	.datab(temp_imemload_output_27),
	.datac(\temp_ALUop_output~0_combout ),
	.datad(\temp_ALUop_output~10_combout ),
	.cin(gnd),
	.combout(\temp_ALUop_output~11_combout ),
	.cout());
// synopsys translate_off
defparam \temp_ALUop_output~11 .lut_mask = 16'hE0A0;
defparam \temp_ALUop_output~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N12
cycloneive_lcell_comb \temp_request_dmemREN_output~0 (
// Equation(s):
// \temp_request_dmemREN_output~0_combout  = (temp_imemload_output_27 & (\temp_branch_output~1_combout  & (temp_imemload_output_26 & !temp_imemload_output_28)))

	.dataa(temp_imemload_output_27),
	.datab(\temp_branch_output~1_combout ),
	.datac(temp_imemload_output_26),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(\temp_request_dmemREN_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_request_dmemREN_output~0 .lut_mask = 16'h0080;
defparam \temp_request_dmemREN_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N20
cycloneive_lcell_comb \temp_request_dmemREN_output~1 (
// Equation(s):
// \temp_request_dmemREN_output~1_combout  = (temp_imemload_output_31 & (!temp_imemload_output_29 & \temp_request_dmemREN_output~0_combout ))

	.dataa(gnd),
	.datab(temp_imemload_output_31),
	.datac(temp_imemload_output_29),
	.datad(\temp_request_dmemREN_output~0_combout ),
	.cin(gnd),
	.combout(\temp_request_dmemREN_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_request_dmemREN_output~1 .lut_mask = 16'h0C00;
defparam \temp_request_dmemREN_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N18
cycloneive_lcell_comb \temp_request_dmemWEN_output~0 (
// Equation(s):
// \temp_request_dmemWEN_output~0_combout  = (temp_imemload_output_31 & (temp_imemload_output_29 & \temp_request_dmemREN_output~0_combout ))

	.dataa(gnd),
	.datab(temp_imemload_output_31),
	.datac(temp_imemload_output_29),
	.datad(\temp_request_dmemREN_output~0_combout ),
	.cin(gnd),
	.combout(\temp_request_dmemWEN_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_request_dmemWEN_output~0 .lut_mask = 16'hC000;
defparam \temp_request_dmemWEN_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N22
cycloneive_lcell_comb \temp_regdst_output~0 (
// Equation(s):
// \temp_regdst_output~0_combout  = (\temp_ALUsrc_output~0_combout  & ((Equal31) # ((temp_imemload_output_5 & WideOr3))))

	.dataa(Equal31),
	.datab(temp_imemload_output_51),
	.datac(\temp_ALUsrc_output~0_combout ),
	.datad(WideOr3),
	.cin(gnd),
	.combout(\temp_regdst_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_regdst_output~0 .lut_mask = 16'hE0A0;
defparam \temp_regdst_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N22
cycloneive_lcell_comb \temp_regwrite_output~0 (
// Equation(s):
// \temp_regwrite_output~0_combout  = (temp_ALUsrc_output & (((!temp_imemload_output_31 & WideOr10)) # (!temp_imemload_output_29))) # (!temp_ALUsrc_output & (!temp_imemload_output_31 & ((WideOr10))))

	.dataa(temp_ALUsrc_output),
	.datab(temp_imemload_output_31),
	.datac(temp_imemload_output_29),
	.datad(WideOr10),
	.cin(gnd),
	.combout(\temp_regwrite_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_regwrite_output~0 .lut_mask = 16'h3B0A;
defparam \temp_regwrite_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N0
cycloneive_lcell_comb \temp_regwrite_output~1 (
// Equation(s):
// \temp_regwrite_output~1_combout  = (\temp_ALUop_output~0_combout  & ((\temp_regdst_output~0_combout ) # ((extended_imm_16 & \temp_regwrite_output~0_combout ))))

	.dataa(extended_imm_16),
	.datab(\temp_regdst_output~0_combout ),
	.datac(\temp_ALUop_output~0_combout ),
	.datad(\temp_regwrite_output~0_combout ),
	.cin(gnd),
	.combout(\temp_regwrite_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_regwrite_output~1 .lut_mask = 16'hE0C0;
defparam \temp_regwrite_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N28
cycloneive_lcell_comb \temp_regdst_output~1 (
// Equation(s):
// \temp_regdst_output~1_combout  = (!temp_imemload_output_31 & (!temp_imemload_output_29 & \temp_request_dmemREN_output~0_combout ))

	.dataa(gnd),
	.datab(temp_imemload_output_31),
	.datac(temp_imemload_output_29),
	.datad(\temp_request_dmemREN_output~0_combout ),
	.cin(gnd),
	.combout(\temp_regdst_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_regdst_output~1 .lut_mask = 16'h0300;
defparam \temp_regdst_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N10
cycloneive_lcell_comb \temp_regdst_output~2 (
// Equation(s):
// \temp_regdst_output~2_combout  = (!id_ex_flush1 & \temp_regdst_output~0_combout )

	.dataa(id_ex_flush),
	.datab(gnd),
	.datac(gnd),
	.datad(\temp_regdst_output~0_combout ),
	.cin(gnd),
	.combout(\temp_regdst_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_regdst_output~2 .lut_mask = 16'h5500;
defparam \temp_regdst_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N10
cycloneive_lcell_comb \temp_request_dmemREN_output~2 (
// Equation(s):
// \temp_request_dmemREN_output~2_combout  = (!temp_imemload_output_29 & \temp_request_dmemREN_output~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(temp_imemload_output_29),
	.datad(\temp_request_dmemREN_output~0_combout ),
	.cin(gnd),
	.combout(\temp_request_dmemREN_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_request_dmemREN_output~2 .lut_mask = 16'h0F00;
defparam \temp_request_dmemREN_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N26
cycloneive_lcell_comb \temp_memtoreg_output~0 (
// Equation(s):
// \temp_memtoreg_output~0_combout  = (!temp_imemload_output_30 & (!temp_imemload_output_31 & (memtoreg & !\temp_ALUsrc_output[0]~2_combout )))

	.dataa(temp_imemload_output_30),
	.datab(temp_imemload_output_31),
	.datac(memtoreg),
	.datad(\temp_ALUsrc_output[0]~2_combout ),
	.cin(gnd),
	.combout(\temp_memtoreg_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_memtoreg_output~0 .lut_mask = 16'h0010;
defparam \temp_memtoreg_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N10
cycloneive_lcell_comb \temp_imemload_output~26 (
// Equation(s):
// \temp_imemload_output~26_combout  = (!ex_mem_flush3 & (temp_imemload_output_31 & !use_after_load))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(temp_imemload_output_31),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~26_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~26 .lut_mask = 16'h0050;
defparam \temp_imemload_output~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N2
cycloneive_lcell_comb \temp_imemload_output~27 (
// Equation(s):
// \temp_imemload_output~27_combout  = (!ex_mem_flush3 & (temp_imemload_output_30 & !use_after_load))

	.dataa(ex_mem_flush),
	.datab(temp_imemload_output_30),
	.datac(gnd),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~27_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~27 .lut_mask = 16'h0044;
defparam \temp_imemload_output~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N20
cycloneive_lcell_comb \temp_imemload_output~28 (
// Equation(s):
// \temp_imemload_output~28_combout  = (!ex_mem_flush3 & (temp_imemload_output_29 & !use_after_load))

	.dataa(ex_mem_flush),
	.datab(temp_imemload_output_29),
	.datac(gnd),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~28_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~28 .lut_mask = 16'h0044;
defparam \temp_imemload_output~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N24
cycloneive_lcell_comb \temp_imemload_output~29 (
// Equation(s):
// \temp_imemload_output~29_combout  = (!use_after_load & (!ex_mem_flush3 & temp_imemload_output_27))

	.dataa(gnd),
	.datab(use_after_load),
	.datac(ex_mem_flush),
	.datad(temp_imemload_output_27),
	.cin(gnd),
	.combout(\temp_imemload_output~29_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~29 .lut_mask = 16'h0300;
defparam \temp_imemload_output~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N10
cycloneive_lcell_comb \temp_imemload_output~30 (
// Equation(s):
// \temp_imemload_output~30_combout  = (temp_imemload_output_26 & (!ex_mem_flush3 & !use_after_load))

	.dataa(temp_imemload_output_26),
	.datab(ex_mem_flush),
	.datac(gnd),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~30_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~30 .lut_mask = 16'h0022;
defparam \temp_imemload_output~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N4
cycloneive_lcell_comb \temp_imemload_output~31 (
// Equation(s):
// \temp_imemload_output~31_combout  = (!ex_mem_flush3 & (temp_imemload_output_28 & !use_after_load))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(temp_imemload_output_28),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_imemload_output~31_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~31 .lut_mask = 16'h0030;
defparam \temp_imemload_output~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N0
cycloneive_lcell_comb \temp_branch_output~2 (
// Equation(s):
// \temp_branch_output~2_combout  = (!temp_imemload_output_27 & (!temp_imemload_output_26 & (!temp_imemload_output_29 & temp_imemload_output_28)))

	.dataa(temp_imemload_output_27),
	.datab(temp_imemload_output_26),
	.datac(temp_imemload_output_29),
	.datad(temp_imemload_output_28),
	.cin(gnd),
	.combout(\temp_branch_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_branch_output~2 .lut_mask = 16'h0100;
defparam \temp_branch_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N18
cycloneive_lcell_comb \temp_branch_output~3 (
// Equation(s):
// \temp_branch_output~3_combout  = (!temp_imemload_output_30 & (!temp_imemload_output_31 & (\temp_branch_output~2_combout  & !\temp_ALUsrc_output[0]~2_combout )))

	.dataa(temp_imemload_output_30),
	.datab(temp_imemload_output_31),
	.datac(\temp_branch_output~2_combout ),
	.datad(\temp_ALUsrc_output[0]~2_combout ),
	.cin(gnd),
	.combout(\temp_branch_output~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_branch_output~3 .lut_mask = 16'h0010;
defparam \temp_branch_output~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N2
cycloneive_lcell_comb \temp_NPC_output~0 (
// Equation(s):
// \temp_NPC_output~0_combout  = (!use_after_load & (temp_NPC_output_1 & !ex_mem_flush3))

	.dataa(use_after_load),
	.datab(gnd),
	.datac(temp_NPC_output_110),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~0 .lut_mask = 16'h0050;
defparam \temp_NPC_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N8
cycloneive_lcell_comb \temp_pcselect_output~0 (
// Equation(s):
// \temp_pcselect_output~0_combout  = (WideOr9 & (!\temp_ALUsrc_output[0]~2_combout  & !temp_imemload_output_31))

	.dataa(WideOr9),
	.datab(\temp_ALUsrc_output[0]~2_combout ),
	.datac(gnd),
	.datad(temp_imemload_output_31),
	.cin(gnd),
	.combout(\temp_pcselect_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_pcselect_output~0 .lut_mask = 16'h0022;
defparam \temp_pcselect_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N8
cycloneive_lcell_comb \temp_pcselect_output~1 (
// Equation(s):
// \temp_pcselect_output~1_combout  = (!temp_imemload_output_0 & (!temp_imemload_output_5 & (!temp_imemload_output_2 & temp_imemload_output_3)))

	.dataa(temp_imemload_output_01),
	.datab(temp_imemload_output_51),
	.datac(temp_imemload_output_210),
	.datad(temp_imemload_output_32),
	.cin(gnd),
	.combout(\temp_pcselect_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_pcselect_output~1 .lut_mask = 16'h0100;
defparam \temp_pcselect_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N30
cycloneive_lcell_comb \temp_pcselect_output~2 (
// Equation(s):
// \temp_pcselect_output~2_combout  = (!temp_imemload_output_1 & (\temp_ALUsrc_output~0_combout  & \temp_pcselect_output~1_combout ))

	.dataa(gnd),
	.datab(temp_imemload_output_110),
	.datac(\temp_ALUsrc_output~0_combout ),
	.datad(\temp_pcselect_output~1_combout ),
	.cin(gnd),
	.combout(\temp_pcselect_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_pcselect_output~2 .lut_mask = 16'h3000;
defparam \temp_pcselect_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N24
cycloneive_lcell_comb \temp_pcselect_output~3 (
// Equation(s):
// \temp_pcselect_output~3_combout  = (\temp_ALUop_output~0_combout  & ((\temp_pcselect_output~2_combout ) # ((Equal3 & temp_imemload_output_27))))

	.dataa(\temp_pcselect_output~2_combout ),
	.datab(\temp_ALUop_output~0_combout ),
	.datac(Equal3),
	.datad(temp_imemload_output_27),
	.cin(gnd),
	.combout(\temp_pcselect_output~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_pcselect_output~3 .lut_mask = 16'hC888;
defparam \temp_pcselect_output~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N24
cycloneive_lcell_comb \temp_NPC_output~1 (
// Equation(s):
// \temp_NPC_output~1_combout  = (!use_after_load & (temp_NPC_output_0 & !ex_mem_flush3))

	.dataa(use_after_load),
	.datab(gnd),
	.datac(temp_NPC_output_01),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~1 .lut_mask = 16'h0050;
defparam \temp_NPC_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N10
cycloneive_lcell_comb \temp_NPC_output~2 (
// Equation(s):
// \temp_NPC_output~2_combout  = (!use_after_load & (temp_NPC_output_2 & !ex_mem_flush3))

	.dataa(use_after_load),
	.datab(gnd),
	.datac(temp_NPC_output_210),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~2 .lut_mask = 16'h0050;
defparam \temp_NPC_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N28
cycloneive_lcell_comb \temp_NPC_output~3 (
// Equation(s):
// \temp_NPC_output~3_combout  = (!ex_mem_flush3 & (!use_after_load & temp_NPC_output_3))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(use_after_load),
	.datad(temp_NPC_output_32),
	.cin(gnd),
	.combout(\temp_NPC_output~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~3 .lut_mask = 16'h0300;
defparam \temp_NPC_output~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N24
cycloneive_lcell_comb \temp_NPC_output~4 (
// Equation(s):
// \temp_NPC_output~4_combout  = (!use_after_load & (temp_NPC_output_5 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(use_after_load),
	.datac(temp_NPC_output_51),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~4 .lut_mask = 16'h0030;
defparam \temp_NPC_output~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N20
cycloneive_lcell_comb \temp_NPC_output~5 (
// Equation(s):
// \temp_NPC_output~5_combout  = (!use_after_load & (!ex_mem_flush3 & temp_NPC_output_4))

	.dataa(use_after_load),
	.datab(ex_mem_flush),
	.datac(temp_NPC_output_41),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~5_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~5 .lut_mask = 16'h1010;
defparam \temp_NPC_output~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N12
cycloneive_lcell_comb \temp_NPC_output~6 (
// Equation(s):
// \temp_NPC_output~6_combout  = (!use_after_load & (temp_NPC_output_7 & !ex_mem_flush3))

	.dataa(use_after_load),
	.datab(gnd),
	.datac(temp_NPC_output_71),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~6_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~6 .lut_mask = 16'h0050;
defparam \temp_NPC_output~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N10
cycloneive_lcell_comb \temp_NPC_output~7 (
// Equation(s):
// \temp_NPC_output~7_combout  = (!ex_mem_flush3 & (temp_NPC_output_6 & !use_after_load))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(temp_NPC_output_61),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_NPC_output~7_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~7 .lut_mask = 16'h0030;
defparam \temp_NPC_output~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N28
cycloneive_lcell_comb \temp_NPC_output~8 (
// Equation(s):
// \temp_NPC_output~8_combout  = (temp_NPC_output_9 & (!ex_mem_flush3 & !use_after_load))

	.dataa(temp_NPC_output_91),
	.datab(gnd),
	.datac(ex_mem_flush),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_NPC_output~8_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~8 .lut_mask = 16'h000A;
defparam \temp_NPC_output~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N6
cycloneive_lcell_comb \temp_NPC_output~9 (
// Equation(s):
// \temp_NPC_output~9_combout  = (!use_after_load & (temp_NPC_output_8 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(use_after_load),
	.datac(temp_NPC_output_81),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~9_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~9 .lut_mask = 16'h0030;
defparam \temp_NPC_output~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N2
cycloneive_lcell_comb \temp_NPC_output~10 (
// Equation(s):
// \temp_NPC_output~10_combout  = (!use_after_load & (temp_NPC_output_11 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(use_after_load),
	.datac(temp_NPC_output_111),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~10_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~10 .lut_mask = 16'h0030;
defparam \temp_NPC_output~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N20
cycloneive_lcell_comb \temp_NPC_output~11 (
// Equation(s):
// \temp_NPC_output~11_combout  = (!use_after_load & (temp_NPC_output_10 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(use_after_load),
	.datac(temp_NPC_output_101),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~11_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~11 .lut_mask = 16'h0030;
defparam \temp_NPC_output~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N16
cycloneive_lcell_comb \temp_NPC_output~12 (
// Equation(s):
// \temp_NPC_output~12_combout  = (!ex_mem_flush3 & (temp_NPC_output_13 & !use_after_load))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(temp_NPC_output_131),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_NPC_output~12_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~12 .lut_mask = 16'h0050;
defparam \temp_NPC_output~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N14
cycloneive_lcell_comb \temp_NPC_output~13 (
// Equation(s):
// \temp_NPC_output~13_combout  = (!ex_mem_flush3 & (temp_NPC_output_12 & !use_after_load))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(temp_NPC_output_121),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_NPC_output~13_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~13 .lut_mask = 16'h0050;
defparam \temp_NPC_output~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N10
cycloneive_lcell_comb \temp_NPC_output~14 (
// Equation(s):
// \temp_NPC_output~14_combout  = (!use_after_load & (temp_NPC_output_15 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(use_after_load),
	.datac(temp_NPC_output_151),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~14_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~14 .lut_mask = 16'h0030;
defparam \temp_NPC_output~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N16
cycloneive_lcell_comb \temp_NPC_output~15 (
// Equation(s):
// \temp_NPC_output~15_combout  = (!use_after_load & (temp_NPC_output_14 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(use_after_load),
	.datac(temp_NPC_output_141),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~15_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~15 .lut_mask = 16'h0030;
defparam \temp_NPC_output~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N0
cycloneive_lcell_comb \temp_NPC_output~16 (
// Equation(s):
// \temp_NPC_output~16_combout  = (!use_after_load & (temp_NPC_output_17 & !ex_mem_flush3))

	.dataa(use_after_load),
	.datab(gnd),
	.datac(temp_NPC_output_171),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~16_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~16 .lut_mask = 16'h0050;
defparam \temp_NPC_output~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N0
cycloneive_lcell_comb \temp_NPC_output~17 (
// Equation(s):
// \temp_NPC_output~17_combout  = (!ex_mem_flush3 & (temp_NPC_output_16 & !use_after_load))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(temp_NPC_output_161),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_NPC_output~17_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~17 .lut_mask = 16'h0030;
defparam \temp_NPC_output~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N12
cycloneive_lcell_comb \temp_NPC_output~18 (
// Equation(s):
// \temp_NPC_output~18_combout  = (!use_after_load & (!ex_mem_flush3 & temp_NPC_output_19))

	.dataa(gnd),
	.datab(use_after_load),
	.datac(ex_mem_flush),
	.datad(temp_NPC_output_191),
	.cin(gnd),
	.combout(\temp_NPC_output~18_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~18 .lut_mask = 16'h0300;
defparam \temp_NPC_output~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N18
cycloneive_lcell_comb \temp_NPC_output~19 (
// Equation(s):
// \temp_NPC_output~19_combout  = (temp_NPC_output_18 & (!ex_mem_flush3 & !use_after_load))

	.dataa(temp_NPC_output_181),
	.datab(ex_mem_flush),
	.datac(use_after_load),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~19_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~19 .lut_mask = 16'h0202;
defparam \temp_NPC_output~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N18
cycloneive_lcell_comb \temp_NPC_output~20 (
// Equation(s):
// \temp_NPC_output~20_combout  = (!use_after_load & (temp_NPC_output_20 & !ex_mem_flush3))

	.dataa(use_after_load),
	.datab(gnd),
	.datac(temp_NPC_output_201),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~20_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~20 .lut_mask = 16'h0050;
defparam \temp_NPC_output~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N4
cycloneive_lcell_comb \temp_NPC_output~21 (
// Equation(s):
// \temp_NPC_output~21_combout  = (!ex_mem_flush3 & (temp_NPC_output_21 & !use_after_load))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(temp_NPC_output_211),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_NPC_output~21_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~21 .lut_mask = 16'h0050;
defparam \temp_NPC_output~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N14
cycloneive_lcell_comb \temp_NPC_output[21]~feeder (
// Equation(s):
// \temp_NPC_output[21]~feeder_combout  = \temp_NPC_output~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\temp_NPC_output~21_combout ),
	.cin(gnd),
	.combout(\temp_NPC_output[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output[21]~feeder .lut_mask = 16'hFF00;
defparam \temp_NPC_output[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N30
cycloneive_lcell_comb \temp_NPC_output~22 (
// Equation(s):
// \temp_NPC_output~22_combout  = (temp_NPC_output_23 & (!use_after_load & !ex_mem_flush3))

	.dataa(temp_NPC_output_231),
	.datab(use_after_load),
	.datac(ex_mem_flush),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~22_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~22 .lut_mask = 16'h0202;
defparam \temp_NPC_output~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N14
cycloneive_lcell_comb \temp_NPC_output~23 (
// Equation(s):
// \temp_NPC_output~23_combout  = (!ex_mem_flush3 & (temp_NPC_output_22 & !use_after_load))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(temp_NPC_output_221),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_NPC_output~23_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~23 .lut_mask = 16'h0030;
defparam \temp_NPC_output~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N0
cycloneive_lcell_comb \temp_NPC_output~24 (
// Equation(s):
// \temp_NPC_output~24_combout  = (!ex_mem_flush3 & (!use_after_load & temp_NPC_output_25))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(use_after_load),
	.datad(temp_NPC_output_251),
	.cin(gnd),
	.combout(\temp_NPC_output~24_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~24 .lut_mask = 16'h0500;
defparam \temp_NPC_output~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N20
cycloneive_lcell_comb \temp_NPC_output~25 (
// Equation(s):
// \temp_NPC_output~25_combout  = (!ex_mem_flush3 & (temp_NPC_output_24 & !use_after_load))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(temp_NPC_output_241),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_NPC_output~25_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~25 .lut_mask = 16'h0030;
defparam \temp_NPC_output~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N0
cycloneive_lcell_comb \temp_NPC_output~26 (
// Equation(s):
// \temp_NPC_output~26_combout  = (!use_after_load & (!ex_mem_flush3 & temp_NPC_output_26))

	.dataa(use_after_load),
	.datab(ex_mem_flush),
	.datac(temp_NPC_output_261),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~26_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~26 .lut_mask = 16'h1010;
defparam \temp_NPC_output~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N20
cycloneive_lcell_comb \temp_NPC_output~27 (
// Equation(s):
// \temp_NPC_output~27_combout  = (!use_after_load & (!ex_mem_flush3 & temp_NPC_output_27))

	.dataa(use_after_load),
	.datab(ex_mem_flush),
	.datac(temp_NPC_output_271),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~27_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~27 .lut_mask = 16'h1010;
defparam \temp_NPC_output~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N16
cycloneive_lcell_comb \temp_NPC_output~28 (
// Equation(s):
// \temp_NPC_output~28_combout  = (!use_after_load & (!ex_mem_flush3 & temp_NPC_output_29))

	.dataa(use_after_load),
	.datab(ex_mem_flush),
	.datac(temp_NPC_output_291),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~28_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~28 .lut_mask = 16'h1010;
defparam \temp_NPC_output~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N14
cycloneive_lcell_comb \temp_NPC_output~29 (
// Equation(s):
// \temp_NPC_output~29_combout  = (!use_after_load & (!ex_mem_flush3 & temp_NPC_output_28))

	.dataa(use_after_load),
	.datab(ex_mem_flush),
	.datac(temp_NPC_output_281),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~29_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~29 .lut_mask = 16'h1010;
defparam \temp_NPC_output~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N30
cycloneive_lcell_comb \temp_NPC_output~30 (
// Equation(s):
// \temp_NPC_output~30_combout  = (!ex_mem_flush3 & (temp_NPC_output_31 & !use_after_load))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(temp_NPC_output_311),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_NPC_output~30_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~30 .lut_mask = 16'h0030;
defparam \temp_NPC_output~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N24
cycloneive_lcell_comb \temp_NPC_output~31 (
// Equation(s):
// \temp_NPC_output~31_combout  = (!ex_mem_flush3 & (temp_NPC_output_30 & !use_after_load))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(temp_NPC_output_301),
	.datad(use_after_load),
	.cin(gnd),
	.combout(\temp_NPC_output~31_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~31 .lut_mask = 16'h0030;
defparam \temp_NPC_output~31 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module if_id_latch (
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	ex_mem_flush,
	Mux30,
	ccifiwait_0,
	temp_imemload_output_17,
	temp_imemload_output_16,
	temp_imemload_output_19,
	temp_imemload_output_18,
	temp_imemload_output_20,
	temp_imemload_output_22,
	temp_imemload_output_21,
	temp_imemload_output_24,
	temp_imemload_output_23,
	temp_imemload_output_25,
	Mux31,
	Mux29,
	Mux28,
	Mux26,
	Mux27,
	Mux24,
	Mux25,
	Mux22,
	Mux23,
	Mux20,
	Mux21,
	Mux18,
	Mux19,
	Mux16,
	Mux17,
	Mux14,
	Mux15,
	Mux12,
	Mux13,
	Mux11,
	Mux10,
	Mux8,
	Mux9,
	Mux6,
	Mux7,
	Mux5,
	Mux4,
	Mux2,
	Mux3,
	Mux0,
	Mux1,
	temp_imemload_output_29,
	temp_imemload_output_31,
	temp_imemload_output_30,
	temp_imemload_output_28,
	temp_imemload_output_27,
	temp_imemload_output_26,
	temp_imemload_output_0,
	temp_imemload_output_2,
	temp_imemload_output_3,
	temp_imemload_output_5,
	temp_imemload_output_15,
	temp_imemload_output_14,
	temp_imemload_output_13,
	temp_imemload_output_12,
	temp_imemload_output_11,
	temp_imemload_output_10,
	temp_imemload_output_9,
	temp_imemload_output_8,
	temp_imemload_output_7,
	temp_imemload_output_6,
	temp_imemload_output_1,
	temp_imemload_output_4,
	wen,
	temp_NPC_output_1,
	temp_NPC_output_0,
	temp_NPC_output_2,
	temp_NPC_output_3,
	temp_NPC_output_5,
	temp_NPC_output_4,
	temp_NPC_output_7,
	temp_NPC_output_6,
	temp_NPC_output_9,
	temp_NPC_output_8,
	temp_NPC_output_11,
	temp_NPC_output_10,
	temp_NPC_output_13,
	temp_NPC_output_12,
	temp_NPC_output_15,
	temp_NPC_output_14,
	temp_NPC_output_17,
	temp_NPC_output_16,
	temp_NPC_output_19,
	temp_NPC_output_18,
	temp_NPC_output_20,
	temp_NPC_output_21,
	temp_NPC_output_23,
	temp_NPC_output_22,
	temp_NPC_output_25,
	temp_NPC_output_24,
	temp_NPC_output_26,
	temp_NPC_output_27,
	temp_NPC_output_29,
	temp_NPC_output_28,
	temp_NPC_output_31,
	temp_NPC_output_30,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	ex_mem_flush;
input 	Mux30;
input 	ccifiwait_0;
output 	temp_imemload_output_17;
output 	temp_imemload_output_16;
output 	temp_imemload_output_19;
output 	temp_imemload_output_18;
output 	temp_imemload_output_20;
output 	temp_imemload_output_22;
output 	temp_imemload_output_21;
output 	temp_imemload_output_24;
output 	temp_imemload_output_23;
output 	temp_imemload_output_25;
input 	Mux31;
input 	Mux29;
input 	Mux28;
input 	Mux26;
input 	Mux27;
input 	Mux24;
input 	Mux25;
input 	Mux22;
input 	Mux23;
input 	Mux20;
input 	Mux21;
input 	Mux18;
input 	Mux19;
input 	Mux16;
input 	Mux17;
input 	Mux14;
input 	Mux15;
input 	Mux12;
input 	Mux13;
input 	Mux11;
input 	Mux10;
input 	Mux8;
input 	Mux9;
input 	Mux6;
input 	Mux7;
input 	Mux5;
input 	Mux4;
input 	Mux2;
input 	Mux3;
input 	Mux0;
input 	Mux1;
output 	temp_imemload_output_29;
output 	temp_imemload_output_31;
output 	temp_imemload_output_30;
output 	temp_imemload_output_28;
output 	temp_imemload_output_27;
output 	temp_imemload_output_26;
output 	temp_imemload_output_0;
output 	temp_imemload_output_2;
output 	temp_imemload_output_3;
output 	temp_imemload_output_5;
output 	temp_imemload_output_15;
output 	temp_imemload_output_14;
output 	temp_imemload_output_13;
output 	temp_imemload_output_12;
output 	temp_imemload_output_11;
output 	temp_imemload_output_10;
output 	temp_imemload_output_9;
output 	temp_imemload_output_8;
output 	temp_imemload_output_7;
output 	temp_imemload_output_6;
output 	temp_imemload_output_1;
output 	temp_imemload_output_4;
input 	wen;
output 	temp_NPC_output_1;
output 	temp_NPC_output_0;
output 	temp_NPC_output_2;
output 	temp_NPC_output_3;
output 	temp_NPC_output_5;
output 	temp_NPC_output_4;
output 	temp_NPC_output_7;
output 	temp_NPC_output_6;
output 	temp_NPC_output_9;
output 	temp_NPC_output_8;
output 	temp_NPC_output_11;
output 	temp_NPC_output_10;
output 	temp_NPC_output_13;
output 	temp_NPC_output_12;
output 	temp_NPC_output_15;
output 	temp_NPC_output_14;
output 	temp_NPC_output_17;
output 	temp_NPC_output_16;
output 	temp_NPC_output_19;
output 	temp_NPC_output_18;
output 	temp_NPC_output_20;
output 	temp_NPC_output_21;
output 	temp_NPC_output_23;
output 	temp_NPC_output_22;
output 	temp_NPC_output_25;
output 	temp_NPC_output_24;
output 	temp_NPC_output_26;
output 	temp_NPC_output_27;
output 	temp_NPC_output_29;
output 	temp_NPC_output_28;
output 	temp_NPC_output_31;
output 	temp_NPC_output_30;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \temp_imemload_output~0_combout ;
wire \temp_imemload_output~1_combout ;
wire \temp_imemload_output~2_combout ;
wire \temp_imemload_output~3_combout ;
wire \temp_imemload_output~4_combout ;
wire \temp_imemload_output~5_combout ;
wire \temp_imemload_output~6_combout ;
wire \temp_imemload_output~7_combout ;
wire \temp_imemload_output~8_combout ;
wire \temp_imemload_output~9_combout ;
wire \temp_imemload_output~10_combout ;
wire \temp_imemload_output~11_combout ;
wire \temp_imemload_output~12_combout ;
wire \temp_imemload_output~13_combout ;
wire \temp_imemload_output~14_combout ;
wire \temp_imemload_output~15_combout ;
wire \temp_imemload_output~16_combout ;
wire \temp_imemload_output~17_combout ;
wire \temp_imemload_output~18_combout ;
wire \temp_imemload_output~19_combout ;
wire \temp_imemload_output~20_combout ;
wire \temp_imemload_output~21_combout ;
wire \temp_imemload_output~22_combout ;
wire \temp_imemload_output~23_combout ;
wire \temp_imemload_output~24_combout ;
wire \temp_imemload_output~25_combout ;
wire \temp_imemload_output~26_combout ;
wire \temp_imemload_output~27_combout ;
wire \temp_imemload_output~28_combout ;
wire \temp_imemload_output~29_combout ;
wire \temp_imemload_output~30_combout ;
wire \temp_imemload_output~31_combout ;
wire \temp_NPC_output~0_combout ;
wire \temp_NPC_output~1_combout ;
wire \temp_NPC_output~2_combout ;
wire \temp_NPC_output~3_combout ;
wire \temp_NPC_output~4_combout ;
wire \temp_NPC_output~5_combout ;
wire \temp_NPC_output~6_combout ;
wire \temp_NPC_output~7_combout ;
wire \temp_NPC_output~8_combout ;
wire \temp_NPC_output~9_combout ;
wire \temp_NPC_output~10_combout ;
wire \temp_NPC_output~11_combout ;
wire \temp_NPC_output~12_combout ;
wire \temp_NPC_output~13_combout ;
wire \temp_NPC_output~14_combout ;
wire \temp_NPC_output~15_combout ;
wire \temp_NPC_output~16_combout ;
wire \temp_NPC_output~17_combout ;
wire \temp_NPC_output~18_combout ;
wire \temp_NPC_output~19_combout ;
wire \temp_NPC_output~20_combout ;
wire \temp_NPC_output~21_combout ;
wire \temp_NPC_output~22_combout ;
wire \temp_NPC_output~23_combout ;
wire \temp_NPC_output~24_combout ;
wire \temp_NPC_output~25_combout ;
wire \temp_NPC_output~26_combout ;
wire \temp_NPC_output~27_combout ;
wire \temp_NPC_output~28_combout ;
wire \temp_NPC_output~29_combout ;
wire \temp_NPC_output~30_combout ;
wire \temp_NPC_output~31_combout ;


// Location: FF_X56_Y44_N9
dffeas \temp_imemload_output[17] (
	.clk(CLK),
	.d(\temp_imemload_output~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[17] .is_wysiwyg = "true";
defparam \temp_imemload_output[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N23
dffeas \temp_imemload_output[16] (
	.clk(CLK),
	.d(\temp_imemload_output~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[16] .is_wysiwyg = "true";
defparam \temp_imemload_output[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N11
dffeas \temp_imemload_output[19] (
	.clk(CLK),
	.d(\temp_imemload_output~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[19] .is_wysiwyg = "true";
defparam \temp_imemload_output[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y43_N3
dffeas \temp_imemload_output[18] (
	.clk(CLK),
	.d(\temp_imemload_output~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[18] .is_wysiwyg = "true";
defparam \temp_imemload_output[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N31
dffeas \temp_imemload_output[20] (
	.clk(CLK),
	.d(\temp_imemload_output~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[20] .is_wysiwyg = "true";
defparam \temp_imemload_output[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N21
dffeas \temp_imemload_output[22] (
	.clk(CLK),
	.d(\temp_imemload_output~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[22] .is_wysiwyg = "true";
defparam \temp_imemload_output[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N19
dffeas \temp_imemload_output[21] (
	.clk(CLK),
	.d(\temp_imemload_output~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[21] .is_wysiwyg = "true";
defparam \temp_imemload_output[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y43_N1
dffeas \temp_imemload_output[24] (
	.clk(CLK),
	.d(\temp_imemload_output~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[24] .is_wysiwyg = "true";
defparam \temp_imemload_output[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N9
dffeas \temp_imemload_output[23] (
	.clk(CLK),
	.d(\temp_imemload_output~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[23] .is_wysiwyg = "true";
defparam \temp_imemload_output[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N5
dffeas \temp_imemload_output[25] (
	.clk(CLK),
	.d(\temp_imemload_output~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[25] .is_wysiwyg = "true";
defparam \temp_imemload_output[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N29
dffeas \temp_imemload_output[29] (
	.clk(CLK),
	.d(\temp_imemload_output~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[29] .is_wysiwyg = "true";
defparam \temp_imemload_output[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N25
dffeas \temp_imemload_output[31] (
	.clk(CLK),
	.d(\temp_imemload_output~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[31] .is_wysiwyg = "true";
defparam \temp_imemload_output[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N31
dffeas \temp_imemload_output[30] (
	.clk(CLK),
	.d(\temp_imemload_output~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[30] .is_wysiwyg = "true";
defparam \temp_imemload_output[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N21
dffeas \temp_imemload_output[28] (
	.clk(CLK),
	.d(\temp_imemload_output~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[28] .is_wysiwyg = "true";
defparam \temp_imemload_output[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N13
dffeas \temp_imemload_output[27] (
	.clk(CLK),
	.d(\temp_imemload_output~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[27] .is_wysiwyg = "true";
defparam \temp_imemload_output[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N29
dffeas \temp_imemload_output[26] (
	.clk(CLK),
	.d(\temp_imemload_output~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[26] .is_wysiwyg = "true";
defparam \temp_imemload_output[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N7
dffeas \temp_imemload_output[0] (
	.clk(CLK),
	.d(\temp_imemload_output~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[0] .is_wysiwyg = "true";
defparam \temp_imemload_output[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N5
dffeas \temp_imemload_output[2] (
	.clk(CLK),
	.d(\temp_imemload_output~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[2] .is_wysiwyg = "true";
defparam \temp_imemload_output[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N19
dffeas \temp_imemload_output[3] (
	.clk(CLK),
	.d(\temp_imemload_output~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[3] .is_wysiwyg = "true";
defparam \temp_imemload_output[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N25
dffeas \temp_imemload_output[5] (
	.clk(CLK),
	.d(\temp_imemload_output~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[5] .is_wysiwyg = "true";
defparam \temp_imemload_output[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N9
dffeas \temp_imemload_output[15] (
	.clk(CLK),
	.d(\temp_imemload_output~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[15] .is_wysiwyg = "true";
defparam \temp_imemload_output[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N23
dffeas \temp_imemload_output[14] (
	.clk(CLK),
	.d(\temp_imemload_output~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[14] .is_wysiwyg = "true";
defparam \temp_imemload_output[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N7
dffeas \temp_imemload_output[13] (
	.clk(CLK),
	.d(\temp_imemload_output~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[13] .is_wysiwyg = "true";
defparam \temp_imemload_output[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N21
dffeas \temp_imemload_output[12] (
	.clk(CLK),
	.d(\temp_imemload_output~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[12] .is_wysiwyg = "true";
defparam \temp_imemload_output[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N3
dffeas \temp_imemload_output[11] (
	.clk(CLK),
	.d(\temp_imemload_output~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[11] .is_wysiwyg = "true";
defparam \temp_imemload_output[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N1
dffeas \temp_imemload_output[10] (
	.clk(CLK),
	.d(\temp_imemload_output~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[10] .is_wysiwyg = "true";
defparam \temp_imemload_output[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N29
dffeas \temp_imemload_output[9] (
	.clk(CLK),
	.d(\temp_imemload_output~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[9] .is_wysiwyg = "true";
defparam \temp_imemload_output[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N19
dffeas \temp_imemload_output[8] (
	.clk(CLK),
	.d(\temp_imemload_output~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[8] .is_wysiwyg = "true";
defparam \temp_imemload_output[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N13
dffeas \temp_imemload_output[7] (
	.clk(CLK),
	.d(\temp_imemload_output~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[7] .is_wysiwyg = "true";
defparam \temp_imemload_output[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N23
dffeas \temp_imemload_output[6] (
	.clk(CLK),
	.d(\temp_imemload_output~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[6] .is_wysiwyg = "true";
defparam \temp_imemload_output[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N9
dffeas \temp_imemload_output[1] (
	.clk(CLK),
	.d(\temp_imemload_output~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[1] .is_wysiwyg = "true";
defparam \temp_imemload_output[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N11
dffeas \temp_imemload_output[4] (
	.clk(CLK),
	.d(\temp_imemload_output~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_imemload_output_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_imemload_output[4] .is_wysiwyg = "true";
defparam \temp_imemload_output[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N27
dffeas \temp_NPC_output[1] (
	.clk(CLK),
	.d(\temp_NPC_output~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[1] .is_wysiwyg = "true";
defparam \temp_NPC_output[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N9
dffeas \temp_NPC_output[0] (
	.clk(CLK),
	.d(\temp_NPC_output~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[0] .is_wysiwyg = "true";
defparam \temp_NPC_output[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N23
dffeas \temp_NPC_output[2] (
	.clk(CLK),
	.d(\temp_NPC_output~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[2] .is_wysiwyg = "true";
defparam \temp_NPC_output[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N13
dffeas \temp_NPC_output[3] (
	.clk(CLK),
	.d(\temp_NPC_output~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[3] .is_wysiwyg = "true";
defparam \temp_NPC_output[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N5
dffeas \temp_NPC_output[5] (
	.clk(CLK),
	.d(\temp_NPC_output~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[5] .is_wysiwyg = "true";
defparam \temp_NPC_output[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y44_N27
dffeas \temp_NPC_output[4] (
	.clk(CLK),
	.d(\temp_NPC_output~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[4] .is_wysiwyg = "true";
defparam \temp_NPC_output[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N31
dffeas \temp_NPC_output[7] (
	.clk(CLK),
	.d(\temp_NPC_output~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[7] .is_wysiwyg = "true";
defparam \temp_NPC_output[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N27
dffeas \temp_NPC_output[6] (
	.clk(CLK),
	.d(\temp_NPC_output~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[6] .is_wysiwyg = "true";
defparam \temp_NPC_output[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N27
dffeas \temp_NPC_output[9] (
	.clk(CLK),
	.d(\temp_NPC_output~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[9] .is_wysiwyg = "true";
defparam \temp_NPC_output[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N15
dffeas \temp_NPC_output[8] (
	.clk(CLK),
	.d(\temp_NPC_output~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[8] .is_wysiwyg = "true";
defparam \temp_NPC_output[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N31
dffeas \temp_NPC_output[11] (
	.clk(CLK),
	.d(\temp_NPC_output~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[11] .is_wysiwyg = "true";
defparam \temp_NPC_output[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N5
dffeas \temp_NPC_output[10] (
	.clk(CLK),
	.d(\temp_NPC_output~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[10] .is_wysiwyg = "true";
defparam \temp_NPC_output[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N27
dffeas \temp_NPC_output[13] (
	.clk(CLK),
	.d(\temp_NPC_output~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[13] .is_wysiwyg = "true";
defparam \temp_NPC_output[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N31
dffeas \temp_NPC_output[12] (
	.clk(CLK),
	.d(\temp_NPC_output~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[12] .is_wysiwyg = "true";
defparam \temp_NPC_output[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N27
dffeas \temp_NPC_output[15] (
	.clk(CLK),
	.d(\temp_NPC_output~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[15] .is_wysiwyg = "true";
defparam \temp_NPC_output[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N9
dffeas \temp_NPC_output[14] (
	.clk(CLK),
	.d(\temp_NPC_output~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[14] .is_wysiwyg = "true";
defparam \temp_NPC_output[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N5
dffeas \temp_NPC_output[17] (
	.clk(CLK),
	.d(\temp_NPC_output~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[17] .is_wysiwyg = "true";
defparam \temp_NPC_output[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N9
dffeas \temp_NPC_output[16] (
	.clk(CLK),
	.d(\temp_NPC_output~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[16] .is_wysiwyg = "true";
defparam \temp_NPC_output[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N5
dffeas \temp_NPC_output[19] (
	.clk(CLK),
	.d(\temp_NPC_output~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[19] .is_wysiwyg = "true";
defparam \temp_NPC_output[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N31
dffeas \temp_NPC_output[18] (
	.clk(CLK),
	.d(\temp_NPC_output~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[18] .is_wysiwyg = "true";
defparam \temp_NPC_output[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N27
dffeas \temp_NPC_output[20] (
	.clk(CLK),
	.d(\temp_NPC_output~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[20] .is_wysiwyg = "true";
defparam \temp_NPC_output[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N23
dffeas \temp_NPC_output[21] (
	.clk(CLK),
	.d(\temp_NPC_output~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[21] .is_wysiwyg = "true";
defparam \temp_NPC_output[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N27
dffeas \temp_NPC_output[23] (
	.clk(CLK),
	.d(\temp_NPC_output~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[23] .is_wysiwyg = "true";
defparam \temp_NPC_output[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y44_N23
dffeas \temp_NPC_output[22] (
	.clk(CLK),
	.d(\temp_NPC_output~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[22] .is_wysiwyg = "true";
defparam \temp_NPC_output[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N7
dffeas \temp_NPC_output[25] (
	.clk(CLK),
	.d(\temp_NPC_output~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[25] .is_wysiwyg = "true";
defparam \temp_NPC_output[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y44_N9
dffeas \temp_NPC_output[24] (
	.clk(CLK),
	.d(\temp_NPC_output~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[24] .is_wysiwyg = "true";
defparam \temp_NPC_output[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N9
dffeas \temp_NPC_output[26] (
	.clk(CLK),
	.d(\temp_NPC_output~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[26] .is_wysiwyg = "true";
defparam \temp_NPC_output[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N27
dffeas \temp_NPC_output[27] (
	.clk(CLK),
	.d(\temp_NPC_output~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[27] .is_wysiwyg = "true";
defparam \temp_NPC_output[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N23
dffeas \temp_NPC_output[29] (
	.clk(CLK),
	.d(\temp_NPC_output~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[29] .is_wysiwyg = "true";
defparam \temp_NPC_output[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N31
dffeas \temp_NPC_output[28] (
	.clk(CLK),
	.d(\temp_NPC_output~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[28] .is_wysiwyg = "true";
defparam \temp_NPC_output[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N23
dffeas \temp_NPC_output[31] (
	.clk(CLK),
	.d(\temp_NPC_output~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[31] .is_wysiwyg = "true";
defparam \temp_NPC_output[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N5
dffeas \temp_NPC_output[30] (
	.clk(CLK),
	.d(\temp_NPC_output~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_NPC_output_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_NPC_output[30] .is_wysiwyg = "true";
defparam \temp_NPC_output[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N8
cycloneive_lcell_comb \temp_imemload_output~0 (
// Equation(s):
// \temp_imemload_output~0_combout  = (!ex_mem_flush3 & (ramiframload_17 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(ramiframload_17),
	.datac(gnd),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~0 .lut_mask = 16'h0044;
defparam \temp_imemload_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N22
cycloneive_lcell_comb \temp_imemload_output~1 (
// Equation(s):
// \temp_imemload_output~1_combout  = (ramiframload_16 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(ramiframload_16),
	.datab(gnd),
	.datac(ex_mem_flush),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~1 .lut_mask = 16'h000A;
defparam \temp_imemload_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N10
cycloneive_lcell_comb \temp_imemload_output~2 (
// Equation(s):
// \temp_imemload_output~2_combout  = (ramiframload_19 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(ramiframload_19),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_imemload_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~2 .lut_mask = 16'h0202;
defparam \temp_imemload_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N2
cycloneive_lcell_comb \temp_imemload_output~3 (
// Equation(s):
// \temp_imemload_output~3_combout  = (!ex_mem_flush3 & (ramiframload_18 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(ramiframload_18),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~3 .lut_mask = 16'h0050;
defparam \temp_imemload_output~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N30
cycloneive_lcell_comb \temp_imemload_output~4 (
// Equation(s):
// \temp_imemload_output~4_combout  = (!ex_mem_flush3 & (ramiframload_20 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(ramiframload_20),
	.datac(gnd),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~4 .lut_mask = 16'h0044;
defparam \temp_imemload_output~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N20
cycloneive_lcell_comb \temp_imemload_output~5 (
// Equation(s):
// \temp_imemload_output~5_combout  = (ramiframload_22 & (!ccifiwait_0 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(ramiframload_22),
	.datac(ccifiwait_0),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_imemload_output~5_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~5 .lut_mask = 16'h000C;
defparam \temp_imemload_output~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N18
cycloneive_lcell_comb \temp_imemload_output~6 (
// Equation(s):
// \temp_imemload_output~6_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & ramiframload_21))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(ccifiwait_0),
	.datad(ramiframload_21),
	.cin(gnd),
	.combout(\temp_imemload_output~6_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~6 .lut_mask = 16'h0500;
defparam \temp_imemload_output~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N0
cycloneive_lcell_comb \temp_imemload_output~7 (
// Equation(s):
// \temp_imemload_output~7_combout  = (ramiframload_24 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(ramiframload_24),
	.datab(ex_mem_flush),
	.datac(gnd),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~7_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~7 .lut_mask = 16'h0022;
defparam \temp_imemload_output~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N8
cycloneive_lcell_comb \temp_imemload_output~8 (
// Equation(s):
// \temp_imemload_output~8_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & ramiframload_23))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(ccifiwait_0),
	.datad(ramiframload_23),
	.cin(gnd),
	.combout(\temp_imemload_output~8_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~8 .lut_mask = 16'h0500;
defparam \temp_imemload_output~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N4
cycloneive_lcell_comb \temp_imemload_output~9 (
// Equation(s):
// \temp_imemload_output~9_combout  = (!ex_mem_flush3 & (ramiframload_25 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(ramiframload_25),
	.datac(ccifiwait_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_imemload_output~9_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~9 .lut_mask = 16'h0404;
defparam \temp_imemload_output~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N28
cycloneive_lcell_comb \temp_imemload_output~10 (
// Equation(s):
// \temp_imemload_output~10_combout  = (!ccifiwait_0 & (!ex_mem_flush3 & ramiframload_29))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(ex_mem_flush),
	.datad(ramiframload_29),
	.cin(gnd),
	.combout(\temp_imemload_output~10_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~10 .lut_mask = 16'h0300;
defparam \temp_imemload_output~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N24
cycloneive_lcell_comb \temp_imemload_output~11 (
// Equation(s):
// \temp_imemload_output~11_combout  = (!ex_mem_flush3 & (ramiframload_31 & !ccifiwait_0))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ramiframload_31),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~11_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~11 .lut_mask = 16'h0030;
defparam \temp_imemload_output~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N30
cycloneive_lcell_comb \temp_imemload_output~12 (
// Equation(s):
// \temp_imemload_output~12_combout  = (ramiframload_30 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(gnd),
	.datab(ramiframload_30),
	.datac(ex_mem_flush),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~12_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~12 .lut_mask = 16'h000C;
defparam \temp_imemload_output~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N20
cycloneive_lcell_comb \temp_imemload_output~13 (
// Equation(s):
// \temp_imemload_output~13_combout  = (ramiframload_28 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(ramiframload_28),
	.datab(ex_mem_flush),
	.datac(gnd),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~13_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~13 .lut_mask = 16'h0022;
defparam \temp_imemload_output~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N12
cycloneive_lcell_comb \temp_imemload_output~14 (
// Equation(s):
// \temp_imemload_output~14_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & ramiframload_27))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(ccifiwait_0),
	.datad(ramiframload_27),
	.cin(gnd),
	.combout(\temp_imemload_output~14_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~14 .lut_mask = 16'h0500;
defparam \temp_imemload_output~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N28
cycloneive_lcell_comb \temp_imemload_output~15 (
// Equation(s):
// \temp_imemload_output~15_combout  = (!ccifiwait_0 & (!ex_mem_flush3 & ramiframload_26))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(ex_mem_flush),
	.datad(ramiframload_26),
	.cin(gnd),
	.combout(\temp_imemload_output~15_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~15 .lut_mask = 16'h0500;
defparam \temp_imemload_output~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N6
cycloneive_lcell_comb \temp_imemload_output~16 (
// Equation(s):
// \temp_imemload_output~16_combout  = (!ccifiwait_0 & (!ex_mem_flush3 & ramiframload_0))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(ex_mem_flush),
	.datad(ramiframload_0),
	.cin(gnd),
	.combout(\temp_imemload_output~16_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~16 .lut_mask = 16'h0500;
defparam \temp_imemload_output~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N4
cycloneive_lcell_comb \temp_imemload_output~17 (
// Equation(s):
// \temp_imemload_output~17_combout  = (!ex_mem_flush3 & (ramiframload_2 & !ccifiwait_0))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ramiframload_2),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~17_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~17 .lut_mask = 16'h0030;
defparam \temp_imemload_output~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N18
cycloneive_lcell_comb \temp_imemload_output~18 (
// Equation(s):
// \temp_imemload_output~18_combout  = (!ex_mem_flush3 & (ramiframload_3 & !ccifiwait_0))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ramiframload_3),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~18_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~18 .lut_mask = 16'h0030;
defparam \temp_imemload_output~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N24
cycloneive_lcell_comb \temp_imemload_output~19 (
// Equation(s):
// \temp_imemload_output~19_combout  = (!ex_mem_flush3 & (ramiframload_5 & !ccifiwait_0))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ramiframload_5),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~19_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~19 .lut_mask = 16'h0030;
defparam \temp_imemload_output~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N8
cycloneive_lcell_comb \temp_imemload_output~20 (
// Equation(s):
// \temp_imemload_output~20_combout  = (ramiframload_15 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(ramiframload_15),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_imemload_output~20_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~20 .lut_mask = 16'h0202;
defparam \temp_imemload_output~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N22
cycloneive_lcell_comb \temp_imemload_output~21 (
// Equation(s):
// \temp_imemload_output~21_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & ramiframload_14))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(ramiframload_14),
	.cin(gnd),
	.combout(\temp_imemload_output~21_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~21 .lut_mask = 16'h0300;
defparam \temp_imemload_output~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N6
cycloneive_lcell_comb \temp_imemload_output~22 (
// Equation(s):
// \temp_imemload_output~22_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & ramiframload_13))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(ramiframload_13),
	.cin(gnd),
	.combout(\temp_imemload_output~22_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~22 .lut_mask = 16'h0300;
defparam \temp_imemload_output~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N20
cycloneive_lcell_comb \temp_imemload_output~23 (
// Equation(s):
// \temp_imemload_output~23_combout  = (ramiframload_12 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(ramiframload_12),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_imemload_output~23_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~23 .lut_mask = 16'h0202;
defparam \temp_imemload_output~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N2
cycloneive_lcell_comb \temp_imemload_output~24 (
// Equation(s):
// \temp_imemload_output~24_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & ramiframload_11))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(ramiframload_11),
	.cin(gnd),
	.combout(\temp_imemload_output~24_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~24 .lut_mask = 16'h0300;
defparam \temp_imemload_output~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N0
cycloneive_lcell_comb \temp_imemload_output~25 (
// Equation(s):
// \temp_imemload_output~25_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & ramiframload_10))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(ramiframload_10),
	.cin(gnd),
	.combout(\temp_imemload_output~25_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~25 .lut_mask = 16'h0300;
defparam \temp_imemload_output~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N28
cycloneive_lcell_comb \temp_imemload_output~26 (
// Equation(s):
// \temp_imemload_output~26_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & ramiframload_9))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(ccifiwait_0),
	.datad(ramiframload_9),
	.cin(gnd),
	.combout(\temp_imemload_output~26_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~26 .lut_mask = 16'h0500;
defparam \temp_imemload_output~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N18
cycloneive_lcell_comb \temp_imemload_output~27 (
// Equation(s):
// \temp_imemload_output~27_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & ramiframload_8))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(ccifiwait_0),
	.datad(ramiframload_8),
	.cin(gnd),
	.combout(\temp_imemload_output~27_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~27 .lut_mask = 16'h0500;
defparam \temp_imemload_output~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N12
cycloneive_lcell_comb \temp_imemload_output~28 (
// Equation(s):
// \temp_imemload_output~28_combout  = (!ex_mem_flush3 & (ramiframload_7 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(ramiframload_7),
	.datac(ccifiwait_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_imemload_output~28_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~28 .lut_mask = 16'h0404;
defparam \temp_imemload_output~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N22
cycloneive_lcell_comb \temp_imemload_output~29 (
// Equation(s):
// \temp_imemload_output~29_combout  = (!ex_mem_flush3 & (ramiframload_6 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(ramiframload_6),
	.datac(ccifiwait_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_imemload_output~29_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~29 .lut_mask = 16'h0404;
defparam \temp_imemload_output~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N8
cycloneive_lcell_comb \temp_imemload_output~30 (
// Equation(s):
// \temp_imemload_output~30_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & ramiframload_1))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(ccifiwait_0),
	.datad(ramiframload_1),
	.cin(gnd),
	.combout(\temp_imemload_output~30_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~30 .lut_mask = 16'h0500;
defparam \temp_imemload_output~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N10
cycloneive_lcell_comb \temp_imemload_output~31 (
// Equation(s):
// \temp_imemload_output~31_combout  = (ramiframload_4 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(ramiframload_4),
	.datab(gnd),
	.datac(ex_mem_flush),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_imemload_output~31_combout ),
	.cout());
// synopsys translate_off
defparam \temp_imemload_output~31 .lut_mask = 16'h000A;
defparam \temp_imemload_output~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N26
cycloneive_lcell_comb \temp_NPC_output~0 (
// Equation(s):
// \temp_NPC_output~0_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux30))

	.dataa(ex_mem_flush),
	.datab(ccifiwait_0),
	.datac(Mux30),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~0 .lut_mask = 16'h1010;
defparam \temp_NPC_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N8
cycloneive_lcell_comb \temp_NPC_output~1 (
// Equation(s):
// \temp_NPC_output~1_combout  = (!ex_mem_flush3 & (Mux31 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(Mux31),
	.datac(ccifiwait_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~1 .lut_mask = 16'h0404;
defparam \temp_NPC_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N22
cycloneive_lcell_comb \temp_NPC_output~2 (
// Equation(s):
// \temp_NPC_output~2_combout  = (!ccifiwait_0 & (Mux29 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(Mux29),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~2 .lut_mask = 16'h0030;
defparam \temp_NPC_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N12
cycloneive_lcell_comb \temp_NPC_output~3 (
// Equation(s):
// \temp_NPC_output~3_combout  = (Mux28 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(Mux28),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~3_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~3 .lut_mask = 16'h0202;
defparam \temp_NPC_output~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N4
cycloneive_lcell_comb \temp_NPC_output~4 (
// Equation(s):
// \temp_NPC_output~4_combout  = (Mux26 & (!ccifiwait_0 & !ex_mem_flush3))

	.dataa(gnd),
	.datab(Mux26),
	.datac(ccifiwait_0),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~4_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~4 .lut_mask = 16'h000C;
defparam \temp_NPC_output~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N26
cycloneive_lcell_comb \temp_NPC_output~5 (
// Equation(s):
// \temp_NPC_output~5_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux27))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux27),
	.cin(gnd),
	.combout(\temp_NPC_output~5_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~5 .lut_mask = 16'h0300;
defparam \temp_NPC_output~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N30
cycloneive_lcell_comb \temp_NPC_output~6 (
// Equation(s):
// \temp_NPC_output~6_combout  = (!ex_mem_flush3 & (Mux24 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(Mux24),
	.datac(ccifiwait_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~6_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~6 .lut_mask = 16'h0404;
defparam \temp_NPC_output~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N26
cycloneive_lcell_comb \temp_NPC_output~7 (
// Equation(s):
// \temp_NPC_output~7_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux25))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux25),
	.cin(gnd),
	.combout(\temp_NPC_output~7_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~7 .lut_mask = 16'h0300;
defparam \temp_NPC_output~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N26
cycloneive_lcell_comb \temp_NPC_output~8 (
// Equation(s):
// \temp_NPC_output~8_combout  = (Mux22 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(Mux22),
	.datab(ex_mem_flush),
	.datac(gnd),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_NPC_output~8_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~8 .lut_mask = 16'h0022;
defparam \temp_NPC_output~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N14
cycloneive_lcell_comb \temp_NPC_output~9 (
// Equation(s):
// \temp_NPC_output~9_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux23))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux23),
	.cin(gnd),
	.combout(\temp_NPC_output~9_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~9 .lut_mask = 16'h0300;
defparam \temp_NPC_output~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N30
cycloneive_lcell_comb \temp_NPC_output~10 (
// Equation(s):
// \temp_NPC_output~10_combout  = (!ccifiwait_0 & (!ex_mem_flush3 & Mux20))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(ex_mem_flush),
	.datad(Mux20),
	.cin(gnd),
	.combout(\temp_NPC_output~10_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~10 .lut_mask = 16'h0500;
defparam \temp_NPC_output~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N4
cycloneive_lcell_comb \temp_NPC_output~11 (
// Equation(s):
// \temp_NPC_output~11_combout  = (!ccifiwait_0 & (Mux21 & !ex_mem_flush3))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(Mux21),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~11_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~11 .lut_mask = 16'h0050;
defparam \temp_NPC_output~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N26
cycloneive_lcell_comb \temp_NPC_output~12 (
// Equation(s):
// \temp_NPC_output~12_combout  = (!ex_mem_flush3 & (Mux18 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(Mux18),
	.datac(gnd),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_NPC_output~12_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~12 .lut_mask = 16'h0044;
defparam \temp_NPC_output~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N30
cycloneive_lcell_comb \temp_NPC_output~13 (
// Equation(s):
// \temp_NPC_output~13_combout  = (!ex_mem_flush3 & (Mux19 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(Mux19),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_NPC_output~13_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~13 .lut_mask = 16'h0050;
defparam \temp_NPC_output~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N26
cycloneive_lcell_comb \temp_NPC_output~14 (
// Equation(s):
// \temp_NPC_output~14_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux16))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux16),
	.cin(gnd),
	.combout(\temp_NPC_output~14_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~14 .lut_mask = 16'h0300;
defparam \temp_NPC_output~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N8
cycloneive_lcell_comb \temp_NPC_output~15 (
// Equation(s):
// \temp_NPC_output~15_combout  = (!ccifiwait_0 & (Mux17 & !ex_mem_flush3))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(Mux17),
	.datad(ex_mem_flush),
	.cin(gnd),
	.combout(\temp_NPC_output~15_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~15 .lut_mask = 16'h0050;
defparam \temp_NPC_output~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N4
cycloneive_lcell_comb \temp_NPC_output~16 (
// Equation(s):
// \temp_NPC_output~16_combout  = (!ex_mem_flush3 & (Mux14 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(Mux14),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_NPC_output~16_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~16 .lut_mask = 16'h0050;
defparam \temp_NPC_output~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N8
cycloneive_lcell_comb \temp_NPC_output~17 (
// Equation(s):
// \temp_NPC_output~17_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux15))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux15),
	.cin(gnd),
	.combout(\temp_NPC_output~17_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~17 .lut_mask = 16'h0300;
defparam \temp_NPC_output~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N4
cycloneive_lcell_comb \temp_NPC_output~18 (
// Equation(s):
// \temp_NPC_output~18_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux12))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux12),
	.cin(gnd),
	.combout(\temp_NPC_output~18_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~18 .lut_mask = 16'h0300;
defparam \temp_NPC_output~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N30
cycloneive_lcell_comb \temp_NPC_output~19 (
// Equation(s):
// \temp_NPC_output~19_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux13))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux13),
	.cin(gnd),
	.combout(\temp_NPC_output~19_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~19 .lut_mask = 16'h0300;
defparam \temp_NPC_output~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N26
cycloneive_lcell_comb \temp_NPC_output~20 (
// Equation(s):
// \temp_NPC_output~20_combout  = (!ex_mem_flush3 & (Mux11 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(Mux11),
	.datac(gnd),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_NPC_output~20_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~20 .lut_mask = 16'h0044;
defparam \temp_NPC_output~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N22
cycloneive_lcell_comb \temp_NPC_output~21 (
// Equation(s):
// \temp_NPC_output~21_combout  = (!ex_mem_flush3 & (Mux10 & !ccifiwait_0))

	.dataa(ex_mem_flush),
	.datab(gnd),
	.datac(Mux10),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_NPC_output~21_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~21 .lut_mask = 16'h0050;
defparam \temp_NPC_output~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N26
cycloneive_lcell_comb \temp_NPC_output~22 (
// Equation(s):
// \temp_NPC_output~22_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux8))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux8),
	.cin(gnd),
	.combout(\temp_NPC_output~22_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~22 .lut_mask = 16'h0300;
defparam \temp_NPC_output~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N22
cycloneive_lcell_comb \temp_NPC_output~23 (
// Equation(s):
// \temp_NPC_output~23_combout  = (Mux9 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(Mux9),
	.datab(ex_mem_flush),
	.datac(gnd),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\temp_NPC_output~23_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~23 .lut_mask = 16'h0022;
defparam \temp_NPC_output~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N6
cycloneive_lcell_comb \temp_NPC_output~24 (
// Equation(s):
// \temp_NPC_output~24_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux6))

	.dataa(ex_mem_flush),
	.datab(ccifiwait_0),
	.datac(Mux6),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~24_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~24 .lut_mask = 16'h1010;
defparam \temp_NPC_output~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N8
cycloneive_lcell_comb \temp_NPC_output~25 (
// Equation(s):
// \temp_NPC_output~25_combout  = (!ccifiwait_0 & (!ex_mem_flush3 & Mux7))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(ex_mem_flush),
	.datad(Mux7),
	.cin(gnd),
	.combout(\temp_NPC_output~25_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~25 .lut_mask = 16'h0300;
defparam \temp_NPC_output~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N8
cycloneive_lcell_comb \temp_NPC_output~26 (
// Equation(s):
// \temp_NPC_output~26_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux5))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux5),
	.cin(gnd),
	.combout(\temp_NPC_output~26_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~26 .lut_mask = 16'h0300;
defparam \temp_NPC_output~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N26
cycloneive_lcell_comb \temp_NPC_output~27 (
// Equation(s):
// \temp_NPC_output~27_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux4))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux4),
	.cin(gnd),
	.combout(\temp_NPC_output~27_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~27 .lut_mask = 16'h0300;
defparam \temp_NPC_output~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N22
cycloneive_lcell_comb \temp_NPC_output~28 (
// Equation(s):
// \temp_NPC_output~28_combout  = (Mux2 & (!ex_mem_flush3 & !ccifiwait_0))

	.dataa(Mux2),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_NPC_output~28_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~28 .lut_mask = 16'h0202;
defparam \temp_NPC_output~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N30
cycloneive_lcell_comb \temp_NPC_output~29 (
// Equation(s):
// \temp_NPC_output~29_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux3))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux3),
	.cin(gnd),
	.combout(\temp_NPC_output~29_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~29 .lut_mask = 16'h0300;
defparam \temp_NPC_output~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N22
cycloneive_lcell_comb \temp_NPC_output~30 (
// Equation(s):
// \temp_NPC_output~30_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux0))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux0),
	.cin(gnd),
	.combout(\temp_NPC_output~30_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~30 .lut_mask = 16'h0300;
defparam \temp_NPC_output~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N4
cycloneive_lcell_comb \temp_NPC_output~31 (
// Equation(s):
// \temp_NPC_output~31_combout  = (!ex_mem_flush3 & (!ccifiwait_0 & Mux1))

	.dataa(gnd),
	.datab(ex_mem_flush),
	.datac(ccifiwait_0),
	.datad(Mux1),
	.cin(gnd),
	.combout(\temp_NPC_output~31_combout ),
	.cout());
// synopsys translate_off
defparam \temp_NPC_output~31 .lut_mask = 16'h0300;
defparam \temp_NPC_output~31 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module mem_to_reg_mux (
	temp_dMemLoad_1,
	temp_aluResult_1,
	temp_memtoreg_0,
	temp_memtoreg_1,
	temp_npc_1,
	Mux30,
	temp_dMemLoad_0,
	temp_aluResult_0,
	temp_npc_0,
	Mux31,
	temp_dMemLoad_2,
	temp_aluResult_2,
	temp_npc_2,
	Mux29,
	temp_dMemLoad_4,
	temp_aluResult_4,
	temp_npc_4,
	Mux27,
	temp_dMemLoad_3,
	temp_aluResult_3,
	temp_npc_3,
	Mux28,
	temp_dMemLoad_8,
	temp_aluResult_8,
	temp_npc_8,
	Mux23,
	temp_dMemLoad_7,
	temp_aluResult_7,
	temp_npc_7,
	Mux24,
	temp_dMemLoad_6,
	temp_aluResult_6,
	temp_npc_6,
	Mux25,
	temp_dMemLoad_5,
	temp_aluResult_5,
	temp_npc_5,
	Mux26,
	temp_dMemLoad_16,
	temp_upper16_16,
	temp_aluResult_16,
	temp_npc_16,
	Mux15,
	temp_dMemLoad_14,
	temp_aluResult_14,
	temp_npc_14,
	Mux17,
	temp_dMemLoad_15,
	temp_aluResult_15,
	temp_npc_15,
	Mux16,
	temp_dMemLoad_13,
	temp_aluResult_13,
	temp_npc_13,
	Mux18,
	temp_dMemLoad_12,
	temp_aluResult_12,
	temp_npc_12,
	Mux19,
	temp_dMemLoad_10,
	temp_aluResult_10,
	temp_npc_10,
	Mux21,
	temp_dMemLoad_11,
	temp_aluResult_11,
	temp_npc_11,
	Mux20,
	temp_dMemLoad_9,
	temp_aluResult_9,
	temp_npc_9,
	Mux22,
	temp_upper16_31,
	temp_dMemLoad_31,
	temp_aluResult_31,
	temp_npc_31,
	Mux0,
	temp_dMemLoad_30,
	temp_upper16_30,
	temp_aluResult_30,
	temp_npc_30,
	Mux1,
	temp_upper16_29,
	temp_dMemLoad_29,
	temp_aluResult_29,
	temp_npc_29,
	Mux2,
	temp_upper16_26,
	temp_dMemLoad_26,
	temp_aluResult_26,
	temp_npc_26,
	Mux5,
	temp_dMemLoad_25,
	temp_upper16_25,
	temp_aluResult_25,
	temp_npc_25,
	Mux6,
	temp_dMemLoad_28,
	temp_upper16_28,
	temp_aluResult_28,
	temp_npc_28,
	Mux3,
	temp_upper16_27,
	temp_dMemLoad_27,
	temp_aluResult_27,
	temp_npc_27,
	Mux4,
	temp_upper16_17,
	temp_dMemLoad_17,
	temp_aluResult_17,
	temp_npc_17,
	Mux14,
	temp_upper16_20,
	temp_dMemLoad_20,
	temp_aluResult_20,
	temp_npc_20,
	Mux11,
	temp_dMemLoad_19,
	temp_upper16_19,
	temp_aluResult_19,
	temp_npc_19,
	Mux12,
	temp_dMemLoad_18,
	temp_upper16_18,
	temp_aluResult_18,
	temp_npc_18,
	Mux13,
	temp_upper16_24,
	temp_dMemLoad_24,
	temp_aluResult_24,
	temp_npc_24,
	Mux7,
	temp_dMemLoad_23,
	temp_upper16_23,
	temp_aluResult_23,
	temp_npc_23,
	Mux8,
	temp_upper16_22,
	temp_dMemLoad_22,
	temp_aluResult_22,
	temp_npc_22,
	Mux9,
	temp_dMemLoad_21,
	temp_upper16_21,
	temp_aluResult_21,
	temp_npc_21,
	Mux10,
	devpor,
	devclrn,
	devoe);
input 	temp_dMemLoad_1;
input 	temp_aluResult_1;
input 	temp_memtoreg_0;
input 	temp_memtoreg_1;
input 	temp_npc_1;
output 	Mux30;
input 	temp_dMemLoad_0;
input 	temp_aluResult_0;
input 	temp_npc_0;
output 	Mux31;
input 	temp_dMemLoad_2;
input 	temp_aluResult_2;
input 	temp_npc_2;
output 	Mux29;
input 	temp_dMemLoad_4;
input 	temp_aluResult_4;
input 	temp_npc_4;
output 	Mux27;
input 	temp_dMemLoad_3;
input 	temp_aluResult_3;
input 	temp_npc_3;
output 	Mux28;
input 	temp_dMemLoad_8;
input 	temp_aluResult_8;
input 	temp_npc_8;
output 	Mux23;
input 	temp_dMemLoad_7;
input 	temp_aluResult_7;
input 	temp_npc_7;
output 	Mux24;
input 	temp_dMemLoad_6;
input 	temp_aluResult_6;
input 	temp_npc_6;
output 	Mux25;
input 	temp_dMemLoad_5;
input 	temp_aluResult_5;
input 	temp_npc_5;
output 	Mux26;
input 	temp_dMemLoad_16;
input 	temp_upper16_16;
input 	temp_aluResult_16;
input 	temp_npc_16;
output 	Mux15;
input 	temp_dMemLoad_14;
input 	temp_aluResult_14;
input 	temp_npc_14;
output 	Mux17;
input 	temp_dMemLoad_15;
input 	temp_aluResult_15;
input 	temp_npc_15;
output 	Mux16;
input 	temp_dMemLoad_13;
input 	temp_aluResult_13;
input 	temp_npc_13;
output 	Mux18;
input 	temp_dMemLoad_12;
input 	temp_aluResult_12;
input 	temp_npc_12;
output 	Mux19;
input 	temp_dMemLoad_10;
input 	temp_aluResult_10;
input 	temp_npc_10;
output 	Mux21;
input 	temp_dMemLoad_11;
input 	temp_aluResult_11;
input 	temp_npc_11;
output 	Mux20;
input 	temp_dMemLoad_9;
input 	temp_aluResult_9;
input 	temp_npc_9;
output 	Mux22;
input 	temp_upper16_31;
input 	temp_dMemLoad_31;
input 	temp_aluResult_31;
input 	temp_npc_31;
output 	Mux0;
input 	temp_dMemLoad_30;
input 	temp_upper16_30;
input 	temp_aluResult_30;
input 	temp_npc_30;
output 	Mux1;
input 	temp_upper16_29;
input 	temp_dMemLoad_29;
input 	temp_aluResult_29;
input 	temp_npc_29;
output 	Mux2;
input 	temp_upper16_26;
input 	temp_dMemLoad_26;
input 	temp_aluResult_26;
input 	temp_npc_26;
output 	Mux5;
input 	temp_dMemLoad_25;
input 	temp_upper16_25;
input 	temp_aluResult_25;
input 	temp_npc_25;
output 	Mux6;
input 	temp_dMemLoad_28;
input 	temp_upper16_28;
input 	temp_aluResult_28;
input 	temp_npc_28;
output 	Mux3;
input 	temp_upper16_27;
input 	temp_dMemLoad_27;
input 	temp_aluResult_27;
input 	temp_npc_27;
output 	Mux4;
input 	temp_upper16_17;
input 	temp_dMemLoad_17;
input 	temp_aluResult_17;
input 	temp_npc_17;
output 	Mux14;
input 	temp_upper16_20;
input 	temp_dMemLoad_20;
input 	temp_aluResult_20;
input 	temp_npc_20;
output 	Mux11;
input 	temp_dMemLoad_19;
input 	temp_upper16_19;
input 	temp_aluResult_19;
input 	temp_npc_19;
output 	Mux12;
input 	temp_dMemLoad_18;
input 	temp_upper16_18;
input 	temp_aluResult_18;
input 	temp_npc_18;
output 	Mux13;
input 	temp_upper16_24;
input 	temp_dMemLoad_24;
input 	temp_aluResult_24;
input 	temp_npc_24;
output 	Mux7;
input 	temp_dMemLoad_23;
input 	temp_upper16_23;
input 	temp_aluResult_23;
input 	temp_npc_23;
output 	Mux8;
input 	temp_upper16_22;
input 	temp_dMemLoad_22;
input 	temp_aluResult_22;
input 	temp_npc_22;
output 	Mux9;
input 	temp_dMemLoad_21;
input 	temp_upper16_21;
input 	temp_aluResult_21;
input 	temp_npc_21;
output 	Mux10;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Mux30~0_combout ;
wire \Mux31~0_combout ;
wire \Mux29~0_combout ;
wire \Mux27~0_combout ;
wire \Mux28~0_combout ;
wire \Mux23~0_combout ;
wire \Mux24~0_combout ;
wire \Mux25~0_combout ;
wire \Mux26~0_combout ;
wire \Mux15~0_combout ;
wire \Mux17~0_combout ;
wire \Mux16~0_combout ;
wire \Mux18~0_combout ;
wire \Mux19~0_combout ;
wire \Mux21~0_combout ;
wire \Mux20~0_combout ;
wire \Mux22~0_combout ;
wire \Mux0~0_combout ;
wire \Mux1~0_combout ;
wire \Mux2~0_combout ;
wire \Mux5~0_combout ;
wire \Mux6~0_combout ;
wire \Mux3~0_combout ;
wire \Mux4~0_combout ;
wire \Mux14~0_combout ;
wire \Mux11~0_combout ;
wire \Mux12~0_combout ;
wire \Mux13~0_combout ;
wire \Mux7~0_combout ;
wire \Mux8~0_combout ;
wire \Mux9~0_combout ;
wire \Mux10~0_combout ;


// Location: LCCOMB_X66_Y44_N24
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// Mux30 = (\Mux30~0_combout ) # ((temp_memtoreg_01 & (temp_memtoreg_11 & temp_npc_1)))

	.dataa(temp_memtoreg_0),
	.datab(temp_memtoreg_1),
	.datac(temp_npc_1),
	.datad(\Mux30~0_combout ),
	.cin(gnd),
	.combout(Mux30),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hFF80;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N28
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// Mux31 = (\Mux31~0_combout ) # ((temp_memtoreg_11 & (temp_memtoreg_01 & temp_npc_0)))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_npc_0),
	.datad(\Mux31~0_combout ),
	.cin(gnd),
	.combout(Mux31),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hFF80;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N16
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// Mux29 = (\Mux29~0_combout ) # ((temp_memtoreg_11 & (temp_npc_2 & temp_memtoreg_01)))

	.dataa(\Mux29~0_combout ),
	.datab(temp_memtoreg_1),
	.datac(temp_npc_2),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(Mux29),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hEAAA;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N12
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// Mux27 = (\Mux27~0_combout ) # ((temp_memtoreg_01 & (temp_memtoreg_11 & temp_npc_4)))

	.dataa(temp_memtoreg_0),
	.datab(\Mux27~0_combout ),
	.datac(temp_memtoreg_1),
	.datad(temp_npc_4),
	.cin(gnd),
	.combout(Mux27),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hECCC;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N16
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// Mux28 = (\Mux28~0_combout ) # ((temp_memtoreg_11 & (temp_npc_3 & temp_memtoreg_01)))

	.dataa(temp_memtoreg_1),
	.datab(temp_npc_3),
	.datac(temp_memtoreg_0),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(Mux28),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hFF80;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N8
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// Mux23 = (\Mux23~0_combout ) # ((temp_npc_8 & (temp_memtoreg_01 & temp_memtoreg_11)))

	.dataa(temp_npc_8),
	.datab(\Mux23~0_combout ),
	.datac(temp_memtoreg_0),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(Mux23),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hECCC;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N12
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// Mux24 = (\Mux24~0_combout ) # ((temp_memtoreg_11 & (temp_npc_7 & temp_memtoreg_01)))

	.dataa(temp_memtoreg_1),
	.datab(\Mux24~0_combout ),
	.datac(temp_npc_7),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(Mux24),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hECCC;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N10
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// Mux25 = (\Mux25~0_combout ) # ((temp_memtoreg_11 & (temp_npc_6 & temp_memtoreg_01)))

	.dataa(temp_memtoreg_1),
	.datab(temp_npc_6),
	.datac(temp_memtoreg_0),
	.datad(\Mux25~0_combout ),
	.cin(gnd),
	.combout(Mux25),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hFF80;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N20
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// Mux26 = (\Mux26~0_combout ) # ((temp_npc_5 & (temp_memtoreg_01 & temp_memtoreg_11)))

	.dataa(temp_npc_5),
	.datab(temp_memtoreg_0),
	.datac(temp_memtoreg_1),
	.datad(\Mux26~0_combout ),
	.cin(gnd),
	.combout(Mux26),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hFF80;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N12
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// Mux15 = (temp_memtoreg_01 & ((\Mux15~0_combout  & ((temp_npc_16))) # (!\Mux15~0_combout  & (temp_dMemLoad_16)))) # (!temp_memtoreg_01 & (((\Mux15~0_combout ))))

	.dataa(temp_dMemLoad_16),
	.datab(temp_npc_16),
	.datac(temp_memtoreg_0),
	.datad(\Mux15~0_combout ),
	.cin(gnd),
	.combout(Mux15),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hCFA0;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N8
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// Mux17 = (\Mux17~0_combout ) # ((temp_npc_14 & (temp_memtoreg_11 & temp_memtoreg_01)))

	.dataa(\Mux17~0_combout ),
	.datab(temp_npc_14),
	.datac(temp_memtoreg_1),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(Mux17),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hEAAA;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N10
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// Mux16 = (\Mux16~0_combout ) # ((temp_npc_15 & (temp_memtoreg_01 & temp_memtoreg_11)))

	.dataa(temp_npc_15),
	.datab(\Mux16~0_combout ),
	.datac(temp_memtoreg_0),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(Mux16),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hECCC;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N30
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// Mux18 = (\Mux18~0_combout ) # ((temp_memtoreg_11 & (temp_npc_13 & temp_memtoreg_01)))

	.dataa(temp_memtoreg_1),
	.datab(temp_npc_13),
	.datac(temp_memtoreg_0),
	.datad(\Mux18~0_combout ),
	.cin(gnd),
	.combout(Mux18),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hFF80;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N24
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// Mux19 = (\Mux19~0_combout ) # ((temp_memtoreg_11 & (temp_memtoreg_01 & temp_npc_12)))

	.dataa(temp_memtoreg_1),
	.datab(\Mux19~0_combout ),
	.datac(temp_memtoreg_0),
	.datad(temp_npc_12),
	.cin(gnd),
	.combout(Mux19),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hECCC;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N28
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// Mux21 = (\Mux21~0_combout ) # ((temp_memtoreg_01 & (temp_memtoreg_11 & temp_npc_10)))

	.dataa(temp_memtoreg_0),
	.datab(temp_memtoreg_1),
	.datac(\Mux21~0_combout ),
	.datad(temp_npc_10),
	.cin(gnd),
	.combout(Mux21),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hF8F0;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N26
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// Mux20 = (\Mux20~0_combout ) # ((temp_memtoreg_11 & (temp_npc_11 & temp_memtoreg_01)))

	.dataa(\Mux20~0_combout ),
	.datab(temp_memtoreg_1),
	.datac(temp_npc_11),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(Mux20),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hEAAA;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N4
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// Mux22 = (\Mux22~0_combout ) # ((temp_npc_9 & (temp_memtoreg_01 & temp_memtoreg_11)))

	.dataa(temp_npc_9),
	.datab(temp_memtoreg_0),
	.datac(temp_memtoreg_1),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(Mux22),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hFF80;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N12
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// Mux0 = (\Mux0~0_combout  & ((temp_npc_31) # ((!temp_memtoreg_11)))) # (!\Mux0~0_combout  & (((temp_memtoreg_11 & temp_upper16_31))))

	.dataa(temp_npc_31),
	.datab(\Mux0~0_combout ),
	.datac(temp_memtoreg_1),
	.datad(temp_upper16_31),
	.cin(gnd),
	.combout(Mux0),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hBC8C;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N12
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// Mux1 = (temp_memtoreg_01 & ((\Mux1~0_combout  & (temp_npc_30)) # (!\Mux1~0_combout  & ((temp_dMemLoad_30))))) # (!temp_memtoreg_01 & (((\Mux1~0_combout ))))

	.dataa(temp_npc_30),
	.datab(temp_memtoreg_0),
	.datac(\Mux1~0_combout ),
	.datad(temp_dMemLoad_30),
	.cin(gnd),
	.combout(Mux1),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hBCB0;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N24
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// Mux2 = (\Mux2~0_combout  & (((temp_npc_29)) # (!temp_memtoreg_11))) # (!\Mux2~0_combout  & (temp_memtoreg_11 & ((temp_upper16_29))))

	.dataa(\Mux2~0_combout ),
	.datab(temp_memtoreg_1),
	.datac(temp_npc_29),
	.datad(temp_upper16_29),
	.cin(gnd),
	.combout(Mux2),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hE6A2;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N8
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// Mux5 = (\Mux5~0_combout  & ((temp_npc_26) # ((!temp_memtoreg_11)))) # (!\Mux5~0_combout  & (((temp_upper16_26 & temp_memtoreg_11))))

	.dataa(\Mux5~0_combout ),
	.datab(temp_npc_26),
	.datac(temp_upper16_26),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(Mux5),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hD8AA;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N6
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// Mux6 = (temp_memtoreg_01 & ((\Mux6~0_combout  & ((temp_npc_25))) # (!\Mux6~0_combout  & (temp_dMemLoad_25)))) # (!temp_memtoreg_01 & (((\Mux6~0_combout ))))

	.dataa(temp_memtoreg_0),
	.datab(temp_dMemLoad_25),
	.datac(temp_npc_25),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(Mux6),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hF588;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N28
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// Mux3 = (temp_memtoreg_01 & ((\Mux3~0_combout  & (temp_npc_28)) # (!\Mux3~0_combout  & ((temp_dMemLoad_28))))) # (!temp_memtoreg_01 & (((\Mux3~0_combout ))))

	.dataa(temp_npc_28),
	.datab(temp_memtoreg_0),
	.datac(temp_dMemLoad_28),
	.datad(\Mux3~0_combout ),
	.cin(gnd),
	.combout(Mux3),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hBBC0;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N26
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// Mux4 = (\Mux4~0_combout  & (((temp_npc_27)) # (!temp_memtoreg_11))) # (!\Mux4~0_combout  & (temp_memtoreg_11 & (temp_upper16_27)))

	.dataa(\Mux4~0_combout ),
	.datab(temp_memtoreg_1),
	.datac(temp_upper16_27),
	.datad(temp_npc_27),
	.cin(gnd),
	.combout(Mux4),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hEA62;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N12
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// Mux14 = (temp_memtoreg_11 & ((\Mux14~0_combout  & (temp_npc_17)) # (!\Mux14~0_combout  & ((temp_upper16_17))))) # (!temp_memtoreg_11 & (((\Mux14~0_combout ))))

	.dataa(temp_memtoreg_1),
	.datab(temp_npc_17),
	.datac(temp_upper16_17),
	.datad(\Mux14~0_combout ),
	.cin(gnd),
	.combout(Mux14),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hDDA0;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N12
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// Mux11 = (temp_memtoreg_11 & ((\Mux11~0_combout  & (temp_npc_20)) # (!\Mux11~0_combout  & ((temp_upper16_20))))) # (!temp_memtoreg_11 & (((\Mux11~0_combout ))))

	.dataa(temp_memtoreg_1),
	.datab(temp_npc_20),
	.datac(temp_upper16_20),
	.datad(\Mux11~0_combout ),
	.cin(gnd),
	.combout(Mux11),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hDDA0;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N14
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// Mux12 = (temp_memtoreg_01 & ((\Mux12~0_combout  & ((temp_npc_19))) # (!\Mux12~0_combout  & (temp_dMemLoad_19)))) # (!temp_memtoreg_01 & (\Mux12~0_combout ))

	.dataa(temp_memtoreg_0),
	.datab(\Mux12~0_combout ),
	.datac(temp_dMemLoad_19),
	.datad(temp_npc_19),
	.cin(gnd),
	.combout(Mux12),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hEC64;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N24
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// Mux13 = (temp_memtoreg_01 & ((\Mux13~0_combout  & (temp_npc_18)) # (!\Mux13~0_combout  & ((temp_dMemLoad_18))))) # (!temp_memtoreg_01 & (((\Mux13~0_combout ))))

	.dataa(temp_npc_18),
	.datab(temp_dMemLoad_18),
	.datac(temp_memtoreg_0),
	.datad(\Mux13~0_combout ),
	.cin(gnd),
	.combout(Mux13),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hAFC0;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N20
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// Mux7 = (temp_memtoreg_11 & ((\Mux7~0_combout  & ((temp_npc_24))) # (!\Mux7~0_combout  & (temp_upper16_24)))) # (!temp_memtoreg_11 & (\Mux7~0_combout ))

	.dataa(temp_memtoreg_1),
	.datab(\Mux7~0_combout ),
	.datac(temp_upper16_24),
	.datad(temp_npc_24),
	.cin(gnd),
	.combout(Mux7),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hEC64;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N16
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// Mux8 = (temp_memtoreg_01 & ((\Mux8~0_combout  & ((temp_npc_23))) # (!\Mux8~0_combout  & (temp_dMemLoad_23)))) # (!temp_memtoreg_01 & (((\Mux8~0_combout ))))

	.dataa(temp_dMemLoad_23),
	.datab(temp_memtoreg_0),
	.datac(\Mux8~0_combout ),
	.datad(temp_npc_23),
	.cin(gnd),
	.combout(Mux8),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hF838;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N22
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// Mux9 = (temp_memtoreg_11 & ((\Mux9~0_combout  & (temp_npc_22)) # (!\Mux9~0_combout  & ((temp_upper16_22))))) # (!temp_memtoreg_11 & (((\Mux9~0_combout ))))

	.dataa(temp_npc_22),
	.datab(temp_memtoreg_1),
	.datac(temp_upper16_22),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(Mux9),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hBBC0;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N8
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// Mux10 = (temp_memtoreg_01 & ((\Mux10~0_combout  & (temp_npc_21)) # (!\Mux10~0_combout  & ((temp_dMemLoad_21))))) # (!temp_memtoreg_01 & (((\Mux10~0_combout ))))

	.dataa(temp_npc_21),
	.datab(temp_memtoreg_0),
	.datac(\Mux10~0_combout ),
	.datad(temp_dMemLoad_21),
	.cin(gnd),
	.combout(Mux10),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hBCB0;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N10
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & ((temp_dMemLoad_1))) # (!temp_memtoreg_01 & (temp_aluResult_110))))

	.dataa(temp_memtoreg_0),
	.datab(temp_memtoreg_1),
	.datac(temp_aluResult_1),
	.datad(temp_dMemLoad_1),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'h3210;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N2
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & ((temp_dMemLoad_0))) # (!temp_memtoreg_01 & (temp_aluResult_01))))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_0),
	.datad(temp_dMemLoad_0),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'h5410;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N22
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_2)) # (!temp_memtoreg_01 & ((temp_aluResult_210)))))

	.dataa(temp_dMemLoad_2),
	.datab(temp_memtoreg_1),
	.datac(temp_aluResult_2),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'h2230;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N0
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_4)) # (!temp_memtoreg_01 & ((temp_aluResult_41)))))

	.dataa(temp_memtoreg_0),
	.datab(temp_dMemLoad_4),
	.datac(temp_aluResult_4),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'h00D8;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N18
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_3)) # (!temp_memtoreg_01 & ((temp_aluResult_32)))))

	.dataa(temp_memtoreg_0),
	.datab(temp_dMemLoad_3),
	.datac(temp_aluResult_3),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'h00D8;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N0
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & ((temp_dMemLoad_8))) # (!temp_memtoreg_01 & (temp_aluResult_81))))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_8),
	.datad(temp_dMemLoad_8),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'h5410;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N2
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_7)) # (!temp_memtoreg_01 & ((temp_aluResult_71)))))

	.dataa(temp_dMemLoad_7),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_7),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'h00B8;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N12
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & ((temp_dMemLoad_6))) # (!temp_memtoreg_01 & (temp_aluResult_61))))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_6),
	.datad(temp_dMemLoad_6),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'h5410;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N18
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & ((temp_dMemLoad_5))) # (!temp_memtoreg_01 & (temp_aluResult_51))))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_5),
	.datad(temp_dMemLoad_5),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'h5410;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N22
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (temp_memtoreg_11 & ((temp_memtoreg_01) # ((temp_upper16_16)))) # (!temp_memtoreg_11 & (!temp_memtoreg_01 & (temp_aluResult_161)))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_16),
	.datad(temp_upper16_16),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hBA98;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N28
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_14)) # (!temp_memtoreg_01 & ((temp_aluResult_141)))))

	.dataa(temp_dMemLoad_14),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_14),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'h00B8;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N0
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_15)) # (!temp_memtoreg_01 & ((temp_aluResult_151)))))

	.dataa(temp_dMemLoad_15),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_15),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'h00B8;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N8
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_13)) # (!temp_memtoreg_01 & ((temp_aluResult_131)))))

	.dataa(temp_memtoreg_0),
	.datab(temp_dMemLoad_13),
	.datac(temp_aluResult_13),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'h00D8;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N6
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_12)) # (!temp_memtoreg_01 & ((temp_aluResult_121)))))

	.dataa(temp_memtoreg_0),
	.datab(temp_dMemLoad_12),
	.datac(temp_aluResult_12),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'h00D8;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N14
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_10)) # (!temp_memtoreg_01 & ((temp_aluResult_101)))))

	.dataa(temp_dMemLoad_10),
	.datab(temp_memtoreg_1),
	.datac(temp_aluResult_10),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'h2230;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N12
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_11)) # (!temp_memtoreg_01 & ((temp_aluResult_111)))))

	.dataa(temp_dMemLoad_11),
	.datab(temp_memtoreg_1),
	.datac(temp_aluResult_11),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'h2230;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N10
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_9)) # (!temp_memtoreg_01 & ((temp_aluResult_91)))))

	.dataa(temp_memtoreg_0),
	.datab(temp_dMemLoad_9),
	.datac(temp_aluResult_9),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'h00D8;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N2
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (temp_memtoreg_01 & ((temp_memtoreg_11) # ((temp_dMemLoad_31)))) # (!temp_memtoreg_01 & (!temp_memtoreg_11 & (temp_aluResult_311)))

	.dataa(temp_memtoreg_0),
	.datab(temp_memtoreg_1),
	.datac(temp_aluResult_31),
	.datad(temp_dMemLoad_31),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hBA98;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N14
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (temp_memtoreg_11 & ((temp_memtoreg_01) # ((temp_upper16_30)))) # (!temp_memtoreg_11 & (!temp_memtoreg_01 & (temp_aluResult_301)))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_30),
	.datad(temp_upper16_30),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hBA98;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N2
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (temp_memtoreg_01 & ((temp_dMemLoad_29) # ((temp_memtoreg_11)))) # (!temp_memtoreg_01 & (((temp_aluResult_291 & !temp_memtoreg_11))))

	.dataa(temp_dMemLoad_29),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_29),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hCCB8;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N10
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (temp_memtoreg_11 & (((temp_memtoreg_01)))) # (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_26)) # (!temp_memtoreg_01 & ((temp_aluResult_261)))))

	.dataa(temp_dMemLoad_26),
	.datab(temp_memtoreg_1),
	.datac(temp_aluResult_26),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hEE30;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N24
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (temp_memtoreg_11 & ((temp_upper16_25) # ((temp_memtoreg_01)))) # (!temp_memtoreg_11 & (((temp_aluResult_251 & !temp_memtoreg_01))))

	.dataa(temp_upper16_25),
	.datab(temp_memtoreg_1),
	.datac(temp_aluResult_25),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hCCB8;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N0
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (temp_memtoreg_01 & (temp_memtoreg_11)) # (!temp_memtoreg_01 & ((temp_memtoreg_11 & ((temp_upper16_28))) # (!temp_memtoreg_11 & (temp_aluResult_281))))

	.dataa(temp_memtoreg_0),
	.datab(temp_memtoreg_1),
	.datac(temp_aluResult_28),
	.datad(temp_upper16_28),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hDC98;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N6
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (temp_memtoreg_11 & (((temp_memtoreg_01)))) # (!temp_memtoreg_11 & ((temp_memtoreg_01 & (temp_dMemLoad_27)) # (!temp_memtoreg_01 & ((temp_aluResult_271)))))

	.dataa(temp_dMemLoad_27),
	.datab(temp_memtoreg_1),
	.datac(temp_aluResult_27),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hEE30;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N22
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (temp_memtoreg_11 & (temp_memtoreg_01)) # (!temp_memtoreg_11 & ((temp_memtoreg_01 & ((temp_dMemLoad_17))) # (!temp_memtoreg_01 & (temp_aluResult_171))))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_17),
	.datad(temp_dMemLoad_17),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hDC98;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N28
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (temp_memtoreg_11 & (temp_memtoreg_01)) # (!temp_memtoreg_11 & ((temp_memtoreg_01 & ((temp_dMemLoad_20))) # (!temp_memtoreg_01 & (temp_aluResult_201))))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_20),
	.datad(temp_dMemLoad_20),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hDC98;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N22
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (temp_memtoreg_11 & ((temp_memtoreg_01) # ((temp_upper16_19)))) # (!temp_memtoreg_11 & (!temp_memtoreg_01 & (temp_aluResult_191)))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_19),
	.datad(temp_upper16_19),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hBA98;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N26
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (temp_memtoreg_11 & ((temp_memtoreg_01) # ((temp_upper16_18)))) # (!temp_memtoreg_11 & (!temp_memtoreg_01 & (temp_aluResult_181)))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_18),
	.datad(temp_upper16_18),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hBA98;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N0
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (temp_memtoreg_11 & (temp_memtoreg_01)) # (!temp_memtoreg_11 & ((temp_memtoreg_01 & ((temp_dMemLoad_24))) # (!temp_memtoreg_01 & (temp_aluResult_241))))

	.dataa(temp_memtoreg_1),
	.datab(temp_memtoreg_0),
	.datac(temp_aluResult_24),
	.datad(temp_dMemLoad_24),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hDC98;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N2
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (temp_memtoreg_01 & (temp_memtoreg_11)) # (!temp_memtoreg_01 & ((temp_memtoreg_11 & ((temp_upper16_23))) # (!temp_memtoreg_11 & (temp_aluResult_231))))

	.dataa(temp_memtoreg_0),
	.datab(temp_memtoreg_1),
	.datac(temp_aluResult_23),
	.datad(temp_upper16_23),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hDC98;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N20
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (temp_memtoreg_01 & ((temp_dMemLoad_22) # ((temp_memtoreg_11)))) # (!temp_memtoreg_01 & (((temp_aluResult_221 & !temp_memtoreg_11))))

	.dataa(temp_memtoreg_0),
	.datab(temp_dMemLoad_22),
	.datac(temp_aluResult_22),
	.datad(temp_memtoreg_1),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hAAD8;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N26
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (temp_memtoreg_01 & (temp_memtoreg_11)) # (!temp_memtoreg_01 & ((temp_memtoreg_11 & ((temp_upper16_21))) # (!temp_memtoreg_11 & (temp_aluResult_211))))

	.dataa(temp_memtoreg_0),
	.datab(temp_memtoreg_1),
	.datac(temp_aluResult_21),
	.datad(temp_upper16_21),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hDC98;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module mem_wb_latch (
	temp_branchDest_0,
	temp_branchDest_4,
	temp_branchDest_3,
	temp_branchDest_2,
	temp_branchDest_1,
	temp_aluResult_1,
	temp_aluResult_0,
	temp_aluResult_2,
	temp_aluResult_3,
	temp_aluResult_5,
	temp_aluResult_4,
	temp_aluResult_7,
	temp_aluResult_6,
	temp_aluResult_9,
	temp_aluResult_8,
	temp_aluResult_11,
	temp_aluResult_10,
	temp_aluResult_13,
	temp_aluResult_12,
	temp_aluResult_15,
	temp_aluResult_14,
	temp_aluResult_17,
	temp_aluResult_16,
	temp_aluResult_19,
	temp_aluResult_18,
	temp_aluResult_20,
	temp_aluResult_21,
	temp_aluResult_23,
	temp_aluResult_22,
	temp_aluResult_25,
	temp_aluResult_24,
	temp_aluResult_26,
	temp_aluResult_27,
	temp_aluResult_29,
	temp_aluResult_28,
	temp_aluResult_31,
	temp_aluResult_30,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	temp_regwrite1,
	temp_memtoreg_0,
	temp_memtoreg_1,
	temp_regwrite2,
	temp_branchDest_11,
	temp_branchDest_01,
	temp_branchDest_31,
	temp_branchDest_21,
	temp_branchDest_41,
	temp_dMemLoad_1,
	temp_aluResult_110,
	temp_memtoreg_01,
	temp_memtoreg_11,
	temp_npc_1,
	temp_dMemLoad_0,
	temp_aluResult_01,
	temp_npc_0,
	temp_dMemLoad_2,
	temp_aluResult_210,
	temp_npc_2,
	temp_dMemLoad_4,
	temp_aluResult_41,
	temp_npc_4,
	temp_dMemLoad_3,
	temp_aluResult_32,
	temp_npc_3,
	temp_dMemLoad_8,
	temp_aluResult_81,
	temp_npc_8,
	temp_dMemLoad_7,
	temp_aluResult_71,
	temp_npc_7,
	temp_dMemLoad_6,
	temp_aluResult_61,
	temp_npc_6,
	temp_dMemLoad_5,
	temp_aluResult_51,
	temp_npc_5,
	temp_dMemLoad_16,
	temp_upper16_16,
	temp_aluResult_161,
	temp_npc_16,
	temp_iMemLoad_0,
	temp_dMemLoad_14,
	temp_aluResult_141,
	temp_npc_14,
	temp_dMemLoad_15,
	temp_aluResult_151,
	temp_npc_15,
	temp_dMemLoad_13,
	temp_aluResult_131,
	temp_npc_13,
	temp_dMemLoad_12,
	temp_aluResult_121,
	temp_npc_12,
	temp_dMemLoad_10,
	temp_aluResult_101,
	temp_npc_10,
	temp_dMemLoad_11,
	temp_aluResult_111,
	temp_npc_11,
	temp_dMemLoad_9,
	temp_aluResult_91,
	temp_npc_9,
	temp_upper16_31,
	temp_dMemLoad_31,
	temp_aluResult_311,
	temp_npc_31,
	temp_iMemLoad_15,
	temp_dMemLoad_30,
	temp_upper16_30,
	temp_aluResult_301,
	temp_npc_30,
	temp_iMemLoad_14,
	temp_upper16_29,
	temp_dMemLoad_29,
	temp_aluResult_291,
	temp_npc_29,
	temp_iMemLoad_13,
	temp_upper16_26,
	temp_dMemLoad_26,
	temp_aluResult_261,
	temp_npc_26,
	temp_iMemLoad_10,
	temp_dMemLoad_25,
	temp_upper16_25,
	temp_aluResult_251,
	temp_npc_25,
	temp_iMemLoad_9,
	temp_dMemLoad_28,
	temp_upper16_28,
	temp_aluResult_281,
	temp_npc_28,
	temp_iMemLoad_12,
	temp_upper16_27,
	temp_dMemLoad_27,
	temp_aluResult_271,
	temp_npc_27,
	temp_iMemLoad_11,
	temp_upper16_17,
	temp_dMemLoad_17,
	temp_aluResult_171,
	temp_npc_17,
	temp_iMemLoad_1,
	temp_upper16_20,
	temp_dMemLoad_20,
	temp_aluResult_201,
	temp_npc_20,
	temp_iMemLoad_4,
	temp_dMemLoad_19,
	temp_upper16_19,
	temp_aluResult_191,
	temp_npc_19,
	temp_iMemLoad_3,
	temp_dMemLoad_18,
	temp_upper16_18,
	temp_aluResult_181,
	temp_npc_18,
	temp_iMemLoad_2,
	temp_upper16_24,
	temp_dMemLoad_24,
	temp_aluResult_241,
	temp_npc_24,
	temp_iMemLoad_8,
	temp_dMemLoad_23,
	temp_upper16_23,
	temp_aluResult_231,
	temp_npc_23,
	temp_iMemLoad_7,
	temp_upper16_22,
	temp_dMemLoad_22,
	temp_aluResult_221,
	temp_npc_22,
	temp_iMemLoad_6,
	temp_dMemLoad_21,
	temp_upper16_21,
	temp_aluResult_211,
	temp_npc_21,
	temp_iMemLoad_5,
	wen,
	temp_npc_110,
	temp_npc_01,
	temp_npc_210,
	temp_npc_32,
	temp_npc_51,
	temp_npc_41,
	temp_npc_71,
	temp_npc_61,
	temp_npc_91,
	temp_npc_81,
	temp_npc_111,
	temp_npc_101,
	temp_npc_131,
	temp_npc_121,
	temp_npc_151,
	temp_npc_141,
	temp_npc_171,
	temp_npc_161,
	temp_npc_191,
	temp_npc_181,
	temp_npc_201,
	temp_npc_211,
	temp_npc_231,
	temp_npc_221,
	temp_npc_251,
	temp_npc_241,
	temp_npc_261,
	temp_npc_271,
	temp_npc_291,
	temp_npc_281,
	temp_npc_311,
	temp_npc_301,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	temp_branchDest_0;
input 	temp_branchDest_4;
input 	temp_branchDest_3;
input 	temp_branchDest_2;
input 	temp_branchDest_1;
input 	temp_aluResult_1;
input 	temp_aluResult_0;
input 	temp_aluResult_2;
input 	temp_aluResult_3;
input 	temp_aluResult_5;
input 	temp_aluResult_4;
input 	temp_aluResult_7;
input 	temp_aluResult_6;
input 	temp_aluResult_9;
input 	temp_aluResult_8;
input 	temp_aluResult_11;
input 	temp_aluResult_10;
input 	temp_aluResult_13;
input 	temp_aluResult_12;
input 	temp_aluResult_15;
input 	temp_aluResult_14;
input 	temp_aluResult_17;
input 	temp_aluResult_16;
input 	temp_aluResult_19;
input 	temp_aluResult_18;
input 	temp_aluResult_20;
input 	temp_aluResult_21;
input 	temp_aluResult_23;
input 	temp_aluResult_22;
input 	temp_aluResult_25;
input 	temp_aluResult_24;
input 	temp_aluResult_26;
input 	temp_aluResult_27;
input 	temp_aluResult_29;
input 	temp_aluResult_28;
input 	temp_aluResult_31;
input 	temp_aluResult_30;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	temp_regwrite1;
input 	temp_memtoreg_0;
input 	temp_memtoreg_1;
output 	temp_regwrite2;
output 	temp_branchDest_11;
output 	temp_branchDest_01;
output 	temp_branchDest_31;
output 	temp_branchDest_21;
output 	temp_branchDest_41;
output 	temp_dMemLoad_1;
output 	temp_aluResult_110;
output 	temp_memtoreg_01;
output 	temp_memtoreg_11;
output 	temp_npc_1;
output 	temp_dMemLoad_0;
output 	temp_aluResult_01;
output 	temp_npc_0;
output 	temp_dMemLoad_2;
output 	temp_aluResult_210;
output 	temp_npc_2;
output 	temp_dMemLoad_4;
output 	temp_aluResult_41;
output 	temp_npc_4;
output 	temp_dMemLoad_3;
output 	temp_aluResult_32;
output 	temp_npc_3;
output 	temp_dMemLoad_8;
output 	temp_aluResult_81;
output 	temp_npc_8;
output 	temp_dMemLoad_7;
output 	temp_aluResult_71;
output 	temp_npc_7;
output 	temp_dMemLoad_6;
output 	temp_aluResult_61;
output 	temp_npc_6;
output 	temp_dMemLoad_5;
output 	temp_aluResult_51;
output 	temp_npc_5;
output 	temp_dMemLoad_16;
output 	temp_upper16_16;
output 	temp_aluResult_161;
output 	temp_npc_16;
input 	temp_iMemLoad_0;
output 	temp_dMemLoad_14;
output 	temp_aluResult_141;
output 	temp_npc_14;
output 	temp_dMemLoad_15;
output 	temp_aluResult_151;
output 	temp_npc_15;
output 	temp_dMemLoad_13;
output 	temp_aluResult_131;
output 	temp_npc_13;
output 	temp_dMemLoad_12;
output 	temp_aluResult_121;
output 	temp_npc_12;
output 	temp_dMemLoad_10;
output 	temp_aluResult_101;
output 	temp_npc_10;
output 	temp_dMemLoad_11;
output 	temp_aluResult_111;
output 	temp_npc_11;
output 	temp_dMemLoad_9;
output 	temp_aluResult_91;
output 	temp_npc_9;
output 	temp_upper16_31;
output 	temp_dMemLoad_31;
output 	temp_aluResult_311;
output 	temp_npc_31;
input 	temp_iMemLoad_15;
output 	temp_dMemLoad_30;
output 	temp_upper16_30;
output 	temp_aluResult_301;
output 	temp_npc_30;
input 	temp_iMemLoad_14;
output 	temp_upper16_29;
output 	temp_dMemLoad_29;
output 	temp_aluResult_291;
output 	temp_npc_29;
input 	temp_iMemLoad_13;
output 	temp_upper16_26;
output 	temp_dMemLoad_26;
output 	temp_aluResult_261;
output 	temp_npc_26;
input 	temp_iMemLoad_10;
output 	temp_dMemLoad_25;
output 	temp_upper16_25;
output 	temp_aluResult_251;
output 	temp_npc_25;
input 	temp_iMemLoad_9;
output 	temp_dMemLoad_28;
output 	temp_upper16_28;
output 	temp_aluResult_281;
output 	temp_npc_28;
input 	temp_iMemLoad_12;
output 	temp_upper16_27;
output 	temp_dMemLoad_27;
output 	temp_aluResult_271;
output 	temp_npc_27;
input 	temp_iMemLoad_11;
output 	temp_upper16_17;
output 	temp_dMemLoad_17;
output 	temp_aluResult_171;
output 	temp_npc_17;
input 	temp_iMemLoad_1;
output 	temp_upper16_20;
output 	temp_dMemLoad_20;
output 	temp_aluResult_201;
output 	temp_npc_20;
input 	temp_iMemLoad_4;
output 	temp_dMemLoad_19;
output 	temp_upper16_19;
output 	temp_aluResult_191;
output 	temp_npc_19;
input 	temp_iMemLoad_3;
output 	temp_dMemLoad_18;
output 	temp_upper16_18;
output 	temp_aluResult_181;
output 	temp_npc_18;
input 	temp_iMemLoad_2;
output 	temp_upper16_24;
output 	temp_dMemLoad_24;
output 	temp_aluResult_241;
output 	temp_npc_24;
input 	temp_iMemLoad_8;
output 	temp_dMemLoad_23;
output 	temp_upper16_23;
output 	temp_aluResult_231;
output 	temp_npc_23;
input 	temp_iMemLoad_7;
output 	temp_upper16_22;
output 	temp_dMemLoad_22;
output 	temp_aluResult_221;
output 	temp_npc_22;
input 	temp_iMemLoad_6;
output 	temp_dMemLoad_21;
output 	temp_upper16_21;
output 	temp_aluResult_211;
output 	temp_npc_21;
input 	temp_iMemLoad_5;
input 	wen;
input 	temp_npc_110;
input 	temp_npc_01;
input 	temp_npc_210;
input 	temp_npc_32;
input 	temp_npc_51;
input 	temp_npc_41;
input 	temp_npc_71;
input 	temp_npc_61;
input 	temp_npc_91;
input 	temp_npc_81;
input 	temp_npc_111;
input 	temp_npc_101;
input 	temp_npc_131;
input 	temp_npc_121;
input 	temp_npc_151;
input 	temp_npc_141;
input 	temp_npc_171;
input 	temp_npc_161;
input 	temp_npc_191;
input 	temp_npc_181;
input 	temp_npc_201;
input 	temp_npc_211;
input 	temp_npc_231;
input 	temp_npc_221;
input 	temp_npc_251;
input 	temp_npc_241;
input 	temp_npc_261;
input 	temp_npc_271;
input 	temp_npc_291;
input 	temp_npc_281;
input 	temp_npc_311;
input 	temp_npc_301;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \temp_dMemLoad[1]~feeder_combout ;
wire \temp_memtoreg[0]~feeder_combout ;
wire \temp_dMemLoad[0]~feeder_combout ;
wire \temp_dMemLoad[2]~feeder_combout ;
wire \temp_dMemLoad[4]~feeder_combout ;
wire \temp_dMemLoad[3]~feeder_combout ;
wire \temp_dMemLoad[8]~feeder_combout ;
wire \temp_npc[8]~feeder_combout ;
wire \temp_npc[7]~feeder_combout ;
wire \temp_dMemLoad[6]~feeder_combout ;
wire \temp_npc[6]~feeder_combout ;
wire \temp_dMemLoad[5]~feeder_combout ;
wire \temp_dMemLoad[16]~feeder_combout ;
wire \temp_upper16[16]~feeder_combout ;
wire \temp_npc[16]~feeder_combout ;
wire \temp_dMemLoad[14]~feeder_combout ;
wire \temp_dMemLoad[15]~feeder_combout ;
wire \temp_npc[15]~feeder_combout ;
wire \temp_dMemLoad[13]~feeder_combout ;
wire \temp_dMemLoad[12]~feeder_combout ;
wire \temp_dMemLoad[10]~feeder_combout ;
wire \temp_npc[10]~feeder_combout ;
wire \temp_dMemLoad[11]~feeder_combout ;
wire \temp_dMemLoad[9]~feeder_combout ;
wire \temp_upper16[31]~feeder_combout ;
wire \temp_dMemLoad[31]~feeder_combout ;
wire \temp_dMemLoad[30]~feeder_combout ;
wire \temp_upper16[30]~feeder_combout ;
wire \temp_upper16[29]~feeder_combout ;
wire \temp_dMemLoad[29]~feeder_combout ;
wire \temp_dMemLoad[26]~feeder_combout ;
wire \temp_dMemLoad[25]~feeder_combout ;
wire \temp_upper16[25]~feeder_combout ;
wire \temp_npc[25]~feeder_combout ;
wire \temp_upper16[28]~feeder_combout ;
wire \temp_dMemLoad[27]~feeder_combout ;
wire \temp_dMemLoad[17]~feeder_combout ;
wire \temp_npc[17]~feeder_combout ;
wire \temp_dMemLoad[20]~feeder_combout ;
wire \temp_npc[20]~feeder_combout ;
wire \temp_upper16[19]~feeder_combout ;
wire \temp_npc[19]~feeder_combout ;
wire \temp_dMemLoad[18]~feeder_combout ;
wire \temp_dMemLoad[24]~feeder_combout ;
wire \temp_dMemLoad[23]~feeder_combout ;
wire \temp_upper16[23]~feeder_combout ;
wire \temp_upper16[22]~feeder_combout ;
wire \temp_dMemLoad[22]~feeder_combout ;
wire \temp_dMemLoad[21]~feeder_combout ;


// Location: FF_X59_Y44_N29
dffeas temp_regwrite(
	.clk(CLK),
	.d(gnd),
	.asdata(temp_regwrite1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_regwrite2),
	.prn(vcc));
// synopsys translate_off
defparam temp_regwrite.is_wysiwyg = "true";
defparam temp_regwrite.power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y44_N9
dffeas \temp_branchDest[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_branchDest_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branchDest_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_branchDest[1] .is_wysiwyg = "true";
defparam \temp_branchDest[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y44_N11
dffeas \temp_branchDest[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_branchDest_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branchDest_01),
	.prn(vcc));
// synopsys translate_off
defparam \temp_branchDest[0] .is_wysiwyg = "true";
defparam \temp_branchDest[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y40_N25
dffeas \temp_branchDest[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_branchDest_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branchDest_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_branchDest[3] .is_wysiwyg = "true";
defparam \temp_branchDest[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N9
dffeas \temp_branchDest[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_branchDest_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branchDest_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_branchDest[2] .is_wysiwyg = "true";
defparam \temp_branchDest[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y40_N13
dffeas \temp_branchDest[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_branchDest_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_branchDest_41),
	.prn(vcc));
// synopsys translate_off
defparam \temp_branchDest[4] .is_wysiwyg = "true";
defparam \temp_branchDest[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y44_N1
dffeas \temp_dMemLoad[1] (
	.clk(CLK),
	.d(\temp_dMemLoad[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[1] .is_wysiwyg = "true";
defparam \temp_dMemLoad[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y44_N11
dffeas \temp_aluResult[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_110),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[1] .is_wysiwyg = "true";
defparam \temp_aluResult[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N9
dffeas \temp_memtoreg[0] (
	.clk(CLK),
	.d(\temp_memtoreg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_memtoreg_01),
	.prn(vcc));
// synopsys translate_off
defparam \temp_memtoreg[0] .is_wysiwyg = "true";
defparam \temp_memtoreg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N13
dffeas \temp_memtoreg[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_memtoreg_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_memtoreg_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_memtoreg[1] .is_wysiwyg = "true";
defparam \temp_memtoreg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y44_N25
dffeas \temp_npc[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_110),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_1),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[1] .is_wysiwyg = "true";
defparam \temp_npc[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N15
dffeas \temp_dMemLoad[0] (
	.clk(CLK),
	.d(\temp_dMemLoad[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[0] .is_wysiwyg = "true";
defparam \temp_dMemLoad[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N3
dffeas \temp_aluResult[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_01),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[0] .is_wysiwyg = "true";
defparam \temp_aluResult[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N29
dffeas \temp_npc[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_01),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_0),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[0] .is_wysiwyg = "true";
defparam \temp_npc[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N5
dffeas \temp_dMemLoad[2] (
	.clk(CLK),
	.d(\temp_dMemLoad[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[2] .is_wysiwyg = "true";
defparam \temp_dMemLoad[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N23
dffeas \temp_aluResult[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_210),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[2] .is_wysiwyg = "true";
defparam \temp_aluResult[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N17
dffeas \temp_npc[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_210),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_2),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[2] .is_wysiwyg = "true";
defparam \temp_npc[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N17
dffeas \temp_dMemLoad[4] (
	.clk(CLK),
	.d(\temp_dMemLoad[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[4] .is_wysiwyg = "true";
defparam \temp_dMemLoad[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N1
dffeas \temp_aluResult[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_41),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[4] .is_wysiwyg = "true";
defparam \temp_aluResult[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y44_N1
dffeas \temp_npc[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_41),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_4),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[4] .is_wysiwyg = "true";
defparam \temp_npc[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N3
dffeas \temp_dMemLoad[3] (
	.clk(CLK),
	.d(\temp_dMemLoad[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[3] .is_wysiwyg = "true";
defparam \temp_dMemLoad[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N19
dffeas \temp_aluResult[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_32),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[3] .is_wysiwyg = "true";
defparam \temp_aluResult[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y37_N9
dffeas \temp_npc[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_32),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_3),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[3] .is_wysiwyg = "true";
defparam \temp_npc[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N7
dffeas \temp_dMemLoad[8] (
	.clk(CLK),
	.d(\temp_dMemLoad[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[8] .is_wysiwyg = "true";
defparam \temp_dMemLoad[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N1
dffeas \temp_aluResult[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_81),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[8] .is_wysiwyg = "true";
defparam \temp_aluResult[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N29
dffeas \temp_npc[8] (
	.clk(CLK),
	.d(\temp_npc[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_8),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[8] .is_wysiwyg = "true";
defparam \temp_npc[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N31
dffeas \temp_dMemLoad[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[7] .is_wysiwyg = "true";
defparam \temp_dMemLoad[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N3
dffeas \temp_aluResult[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_71),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[7] .is_wysiwyg = "true";
defparam \temp_aluResult[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N5
dffeas \temp_npc[7] (
	.clk(CLK),
	.d(\temp_npc[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_7),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[7] .is_wysiwyg = "true";
defparam \temp_npc[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N7
dffeas \temp_dMemLoad[6] (
	.clk(CLK),
	.d(\temp_dMemLoad[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[6] .is_wysiwyg = "true";
defparam \temp_dMemLoad[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N13
dffeas \temp_aluResult[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_61),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[6] .is_wysiwyg = "true";
defparam \temp_aluResult[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N29
dffeas \temp_npc[6] (
	.clk(CLK),
	.d(\temp_npc[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_6),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[6] .is_wysiwyg = "true";
defparam \temp_npc[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N21
dffeas \temp_dMemLoad[5] (
	.clk(CLK),
	.d(\temp_dMemLoad[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[5] .is_wysiwyg = "true";
defparam \temp_dMemLoad[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N19
dffeas \temp_aluResult[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_51),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[5] .is_wysiwyg = "true";
defparam \temp_aluResult[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N27
dffeas \temp_npc[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_51),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_5),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[5] .is_wysiwyg = "true";
defparam \temp_npc[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N31
dffeas \temp_dMemLoad[16] (
	.clk(CLK),
	.d(\temp_dMemLoad[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[16] .is_wysiwyg = "true";
defparam \temp_dMemLoad[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N13
dffeas \temp_upper16[16] (
	.clk(CLK),
	.d(\temp_upper16[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[16] .is_wysiwyg = "true";
defparam \temp_upper16[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N23
dffeas \temp_aluResult[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_161),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[16] .is_wysiwyg = "true";
defparam \temp_aluResult[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y45_N19
dffeas \temp_npc[16] (
	.clk(CLK),
	.d(\temp_npc[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_16),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[16] .is_wysiwyg = "true";
defparam \temp_npc[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N3
dffeas \temp_dMemLoad[14] (
	.clk(CLK),
	.d(\temp_dMemLoad[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[14] .is_wysiwyg = "true";
defparam \temp_dMemLoad[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N29
dffeas \temp_aluResult[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_141),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[14] .is_wysiwyg = "true";
defparam \temp_aluResult[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N13
dffeas \temp_npc[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_141),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_14),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[14] .is_wysiwyg = "true";
defparam \temp_npc[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N7
dffeas \temp_dMemLoad[15] (
	.clk(CLK),
	.d(\temp_dMemLoad[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[15] .is_wysiwyg = "true";
defparam \temp_dMemLoad[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N1
dffeas \temp_aluResult[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_151),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[15] .is_wysiwyg = "true";
defparam \temp_aluResult[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y45_N31
dffeas \temp_npc[15] (
	.clk(CLK),
	.d(\temp_npc[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_15),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[15] .is_wysiwyg = "true";
defparam \temp_npc[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N25
dffeas \temp_dMemLoad[13] (
	.clk(CLK),
	.d(\temp_dMemLoad[13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[13] .is_wysiwyg = "true";
defparam \temp_dMemLoad[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N9
dffeas \temp_aluResult[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_131),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[13] .is_wysiwyg = "true";
defparam \temp_aluResult[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N25
dffeas \temp_npc[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_131),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_13),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[13] .is_wysiwyg = "true";
defparam \temp_npc[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N21
dffeas \temp_dMemLoad[12] (
	.clk(CLK),
	.d(\temp_dMemLoad[12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[12] .is_wysiwyg = "true";
defparam \temp_dMemLoad[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N7
dffeas \temp_aluResult[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_121),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[12] .is_wysiwyg = "true";
defparam \temp_aluResult[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N19
dffeas \temp_npc[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_121),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_12),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[12] .is_wysiwyg = "true";
defparam \temp_npc[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N17
dffeas \temp_dMemLoad[10] (
	.clk(CLK),
	.d(\temp_dMemLoad[10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[10] .is_wysiwyg = "true";
defparam \temp_dMemLoad[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N15
dffeas \temp_aluResult[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_101),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[10] .is_wysiwyg = "true";
defparam \temp_aluResult[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y42_N25
dffeas \temp_npc[10] (
	.clk(CLK),
	.d(\temp_npc[10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_10),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[10] .is_wysiwyg = "true";
defparam \temp_npc[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N31
dffeas \temp_dMemLoad[11] (
	.clk(CLK),
	.d(\temp_dMemLoad[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[11] .is_wysiwyg = "true";
defparam \temp_dMemLoad[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N13
dffeas \temp_aluResult[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_111),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[11] .is_wysiwyg = "true";
defparam \temp_aluResult[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N27
dffeas \temp_npc[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_111),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_11),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[11] .is_wysiwyg = "true";
defparam \temp_npc[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N11
dffeas \temp_dMemLoad[9] (
	.clk(CLK),
	.d(\temp_dMemLoad[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[9] .is_wysiwyg = "true";
defparam \temp_dMemLoad[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N11
dffeas \temp_aluResult[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_91),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[9] .is_wysiwyg = "true";
defparam \temp_aluResult[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N5
dffeas \temp_npc[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_91),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_9),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[9] .is_wysiwyg = "true";
defparam \temp_npc[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N17
dffeas \temp_upper16[31] (
	.clk(CLK),
	.d(\temp_upper16[31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[31] .is_wysiwyg = "true";
defparam \temp_upper16[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N21
dffeas \temp_dMemLoad[31] (
	.clk(CLK),
	.d(\temp_dMemLoad[31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[31] .is_wysiwyg = "true";
defparam \temp_dMemLoad[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N3
dffeas \temp_aluResult[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_311),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[31] .is_wysiwyg = "true";
defparam \temp_aluResult[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y44_N15
dffeas \temp_npc[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_311),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_31),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[31] .is_wysiwyg = "true";
defparam \temp_npc[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N13
dffeas \temp_dMemLoad[30] (
	.clk(CLK),
	.d(\temp_dMemLoad[30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[30] .is_wysiwyg = "true";
defparam \temp_dMemLoad[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N1
dffeas \temp_upper16[30] (
	.clk(CLK),
	.d(\temp_upper16[30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[30] .is_wysiwyg = "true";
defparam \temp_upper16[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N15
dffeas \temp_aluResult[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_301),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[30] .is_wysiwyg = "true";
defparam \temp_aluResult[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y44_N27
dffeas \temp_npc[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_301),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_30),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[30] .is_wysiwyg = "true";
defparam \temp_npc[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N7
dffeas \temp_upper16[29] (
	.clk(CLK),
	.d(\temp_upper16[29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[29] .is_wysiwyg = "true";
defparam \temp_upper16[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N5
dffeas \temp_dMemLoad[29] (
	.clk(CLK),
	.d(\temp_dMemLoad[29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[29] .is_wysiwyg = "true";
defparam \temp_dMemLoad[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N3
dffeas \temp_aluResult[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_291),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[29] .is_wysiwyg = "true";
defparam \temp_aluResult[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N25
dffeas \temp_npc[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_291),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_29),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[29] .is_wysiwyg = "true";
defparam \temp_npc[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N9
dffeas \temp_upper16[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_iMemLoad_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[26] .is_wysiwyg = "true";
defparam \temp_upper16[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N9
dffeas \temp_dMemLoad[26] (
	.clk(CLK),
	.d(\temp_dMemLoad[26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[26] .is_wysiwyg = "true";
defparam \temp_dMemLoad[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N11
dffeas \temp_aluResult[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_261),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[26] .is_wysiwyg = "true";
defparam \temp_aluResult[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N29
dffeas \temp_npc[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_261),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_26),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[26] .is_wysiwyg = "true";
defparam \temp_npc[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N17
dffeas \temp_dMemLoad[25] (
	.clk(CLK),
	.d(\temp_dMemLoad[25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[25] .is_wysiwyg = "true";
defparam \temp_dMemLoad[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N31
dffeas \temp_upper16[25] (
	.clk(CLK),
	.d(\temp_upper16[25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[25] .is_wysiwyg = "true";
defparam \temp_upper16[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N25
dffeas \temp_aluResult[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_251),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[25] .is_wysiwyg = "true";
defparam \temp_aluResult[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N9
dffeas \temp_npc[25] (
	.clk(CLK),
	.d(\temp_npc[25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_25),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[25] .is_wysiwyg = "true";
defparam \temp_npc[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y40_N29
dffeas \temp_dMemLoad[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[28] .is_wysiwyg = "true";
defparam \temp_dMemLoad[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N11
dffeas \temp_upper16[28] (
	.clk(CLK),
	.d(\temp_upper16[28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[28] .is_wysiwyg = "true";
defparam \temp_upper16[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N1
dffeas \temp_aluResult[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_281),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[28] .is_wysiwyg = "true";
defparam \temp_aluResult[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y40_N7
dffeas \temp_npc[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_281),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_28),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[28] .is_wysiwyg = "true";
defparam \temp_npc[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N27
dffeas \temp_upper16[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_iMemLoad_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[27] .is_wysiwyg = "true";
defparam \temp_upper16[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N25
dffeas \temp_dMemLoad[27] (
	.clk(CLK),
	.d(\temp_dMemLoad[27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[27] .is_wysiwyg = "true";
defparam \temp_dMemLoad[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N7
dffeas \temp_aluResult[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_271),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[27] .is_wysiwyg = "true";
defparam \temp_aluResult[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N25
dffeas \temp_npc[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_271),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_27),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[27] .is_wysiwyg = "true";
defparam \temp_npc[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N11
dffeas \temp_upper16[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_iMemLoad_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[17] .is_wysiwyg = "true";
defparam \temp_upper16[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N13
dffeas \temp_dMemLoad[17] (
	.clk(CLK),
	.d(\temp_dMemLoad[17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[17] .is_wysiwyg = "true";
defparam \temp_dMemLoad[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N23
dffeas \temp_aluResult[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_171),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[17] .is_wysiwyg = "true";
defparam \temp_aluResult[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N25
dffeas \temp_npc[17] (
	.clk(CLK),
	.d(\temp_npc[17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_17),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[17] .is_wysiwyg = "true";
defparam \temp_npc[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N13
dffeas \temp_upper16[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_iMemLoad_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[20] .is_wysiwyg = "true";
defparam \temp_upper16[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N11
dffeas \temp_dMemLoad[20] (
	.clk(CLK),
	.d(\temp_dMemLoad[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[20] .is_wysiwyg = "true";
defparam \temp_dMemLoad[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N29
dffeas \temp_aluResult[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_201),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[20] .is_wysiwyg = "true";
defparam \temp_aluResult[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y44_N3
dffeas \temp_npc[20] (
	.clk(CLK),
	.d(\temp_npc[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_20),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[20] .is_wysiwyg = "true";
defparam \temp_npc[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N15
dffeas \temp_dMemLoad[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[19] .is_wysiwyg = "true";
defparam \temp_dMemLoad[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N25
dffeas \temp_upper16[19] (
	.clk(CLK),
	.d(\temp_upper16[19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[19] .is_wysiwyg = "true";
defparam \temp_upper16[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N23
dffeas \temp_aluResult[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_191),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[19] .is_wysiwyg = "true";
defparam \temp_aluResult[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N1
dffeas \temp_npc[19] (
	.clk(CLK),
	.d(\temp_npc[19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_19),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[19] .is_wysiwyg = "true";
defparam \temp_npc[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y43_N29
dffeas \temp_dMemLoad[18] (
	.clk(CLK),
	.d(\temp_dMemLoad[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[18] .is_wysiwyg = "true";
defparam \temp_dMemLoad[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N17
dffeas \temp_upper16[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_iMemLoad_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[18] .is_wysiwyg = "true";
defparam \temp_upper16[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N27
dffeas \temp_aluResult[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_181),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[18] .is_wysiwyg = "true";
defparam \temp_aluResult[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y44_N21
dffeas \temp_npc[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_181),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_18),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[18] .is_wysiwyg = "true";
defparam \temp_npc[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N21
dffeas \temp_upper16[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_iMemLoad_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[24] .is_wysiwyg = "true";
defparam \temp_upper16[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N19
dffeas \temp_dMemLoad[24] (
	.clk(CLK),
	.d(\temp_dMemLoad[24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[24] .is_wysiwyg = "true";
defparam \temp_dMemLoad[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y43_N1
dffeas \temp_aluResult[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_241),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[24] .is_wysiwyg = "true";
defparam \temp_aluResult[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y44_N13
dffeas \temp_npc[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_241),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_24),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[24] .is_wysiwyg = "true";
defparam \temp_npc[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N17
dffeas \temp_dMemLoad[23] (
	.clk(CLK),
	.d(\temp_dMemLoad[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[23] .is_wysiwyg = "true";
defparam \temp_dMemLoad[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N13
dffeas \temp_upper16[23] (
	.clk(CLK),
	.d(\temp_upper16[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[23] .is_wysiwyg = "true";
defparam \temp_upper16[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N3
dffeas \temp_aluResult[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_231),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[23] .is_wysiwyg = "true";
defparam \temp_aluResult[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y44_N31
dffeas \temp_npc[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_231),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_23),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[23] .is_wysiwyg = "true";
defparam \temp_npc[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N15
dffeas \temp_upper16[22] (
	.clk(CLK),
	.d(\temp_upper16[22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[22] .is_wysiwyg = "true";
defparam \temp_upper16[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N19
dffeas \temp_dMemLoad[22] (
	.clk(CLK),
	.d(\temp_dMemLoad[22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[22] .is_wysiwyg = "true";
defparam \temp_dMemLoad[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N21
dffeas \temp_aluResult[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_221),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[22] .is_wysiwyg = "true";
defparam \temp_aluResult[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y44_N9
dffeas \temp_npc[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_221),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_22),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[22] .is_wysiwyg = "true";
defparam \temp_npc[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N15
dffeas \temp_dMemLoad[21] (
	.clk(CLK),
	.d(\temp_dMemLoad[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_dMemLoad_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_dMemLoad[21] .is_wysiwyg = "true";
defparam \temp_dMemLoad[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N1
dffeas \temp_upper16[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_iMemLoad_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_upper16_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_upper16[21] .is_wysiwyg = "true";
defparam \temp_upper16[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y41_N27
dffeas \temp_aluResult[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_aluResult_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_aluResult_211),
	.prn(vcc));
// synopsys translate_off
defparam \temp_aluResult[21] .is_wysiwyg = "true";
defparam \temp_aluResult[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N11
dffeas \temp_npc[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(temp_npc_211),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(temp_npc_21),
	.prn(vcc));
// synopsys translate_off
defparam \temp_npc[21] .is_wysiwyg = "true";
defparam \temp_npc[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y44_N0
cycloneive_lcell_comb \temp_dMemLoad[1]~feeder (
// Equation(s):
// \temp_dMemLoad[1]~feeder_combout  = ramiframload_1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_1),
	.cin(gnd),
	.combout(\temp_dMemLoad[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[1]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N8
cycloneive_lcell_comb \temp_memtoreg[0]~feeder (
// Equation(s):
// \temp_memtoreg[0]~feeder_combout  = temp_memtoreg_0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_memtoreg_0),
	.cin(gnd),
	.combout(\temp_memtoreg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_memtoreg[0]~feeder .lut_mask = 16'hFF00;
defparam \temp_memtoreg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N14
cycloneive_lcell_comb \temp_dMemLoad[0]~feeder (
// Equation(s):
// \temp_dMemLoad[0]~feeder_combout  = ramiframload_0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_0),
	.cin(gnd),
	.combout(\temp_dMemLoad[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[0]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N4
cycloneive_lcell_comb \temp_dMemLoad[2]~feeder (
// Equation(s):
// \temp_dMemLoad[2]~feeder_combout  = ramiframload_2

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_2),
	.cin(gnd),
	.combout(\temp_dMemLoad[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[2]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N16
cycloneive_lcell_comb \temp_dMemLoad[4]~feeder (
// Equation(s):
// \temp_dMemLoad[4]~feeder_combout  = ramiframload_4

	.dataa(ramiframload_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_dMemLoad[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[4]~feeder .lut_mask = 16'hAAAA;
defparam \temp_dMemLoad[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N2
cycloneive_lcell_comb \temp_dMemLoad[3]~feeder (
// Equation(s):
// \temp_dMemLoad[3]~feeder_combout  = ramiframload_3

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_dMemLoad[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[3]~feeder .lut_mask = 16'hF0F0;
defparam \temp_dMemLoad[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N6
cycloneive_lcell_comb \temp_dMemLoad[8]~feeder (
// Equation(s):
// \temp_dMemLoad[8]~feeder_combout  = ramiframload_8

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_8),
	.cin(gnd),
	.combout(\temp_dMemLoad[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[8]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N28
cycloneive_lcell_comb \temp_npc[8]~feeder (
// Equation(s):
// \temp_npc[8]~feeder_combout  = temp_npc_8

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_npc_81),
	.cin(gnd),
	.combout(\temp_npc[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc[8]~feeder .lut_mask = 16'hFF00;
defparam \temp_npc[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N4
cycloneive_lcell_comb \temp_npc[7]~feeder (
// Equation(s):
// \temp_npc[7]~feeder_combout  = temp_npc_7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_npc_71),
	.cin(gnd),
	.combout(\temp_npc[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc[7]~feeder .lut_mask = 16'hFF00;
defparam \temp_npc[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N6
cycloneive_lcell_comb \temp_dMemLoad[6]~feeder (
// Equation(s):
// \temp_dMemLoad[6]~feeder_combout  = ramiframload_6

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_6),
	.cin(gnd),
	.combout(\temp_dMemLoad[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[6]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N28
cycloneive_lcell_comb \temp_npc[6]~feeder (
// Equation(s):
// \temp_npc[6]~feeder_combout  = temp_npc_6

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_npc_61),
	.cin(gnd),
	.combout(\temp_npc[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc[6]~feeder .lut_mask = 16'hFF00;
defparam \temp_npc[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N20
cycloneive_lcell_comb \temp_dMemLoad[5]~feeder (
// Equation(s):
// \temp_dMemLoad[5]~feeder_combout  = ramiframload_5

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_5),
	.cin(gnd),
	.combout(\temp_dMemLoad[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[5]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N30
cycloneive_lcell_comb \temp_dMemLoad[16]~feeder (
// Equation(s):
// \temp_dMemLoad[16]~feeder_combout  = ramiframload_16

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(\temp_dMemLoad[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[16]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N12
cycloneive_lcell_comb \temp_upper16[16]~feeder (
// Equation(s):
// \temp_upper16[16]~feeder_combout  = temp_iMemLoad_0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_iMemLoad_0),
	.cin(gnd),
	.combout(\temp_upper16[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_upper16[16]~feeder .lut_mask = 16'hFF00;
defparam \temp_upper16[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y45_N18
cycloneive_lcell_comb \temp_npc[16]~feeder (
// Equation(s):
// \temp_npc[16]~feeder_combout  = temp_npc_16

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_npc_161),
	.cin(gnd),
	.combout(\temp_npc[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc[16]~feeder .lut_mask = 16'hFF00;
defparam \temp_npc[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N2
cycloneive_lcell_comb \temp_dMemLoad[14]~feeder (
// Equation(s):
// \temp_dMemLoad[14]~feeder_combout  = ramiframload_14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_14),
	.cin(gnd),
	.combout(\temp_dMemLoad[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[14]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N6
cycloneive_lcell_comb \temp_dMemLoad[15]~feeder (
// Equation(s):
// \temp_dMemLoad[15]~feeder_combout  = ramiframload_15

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_15),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_dMemLoad[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[15]~feeder .lut_mask = 16'hF0F0;
defparam \temp_dMemLoad[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y45_N30
cycloneive_lcell_comb \temp_npc[15]~feeder (
// Equation(s):
// \temp_npc[15]~feeder_combout  = temp_npc_15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_npc_151),
	.cin(gnd),
	.combout(\temp_npc[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc[15]~feeder .lut_mask = 16'hFF00;
defparam \temp_npc[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N24
cycloneive_lcell_comb \temp_dMemLoad[13]~feeder (
// Equation(s):
// \temp_dMemLoad[13]~feeder_combout  = ramiframload_13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_13),
	.cin(gnd),
	.combout(\temp_dMemLoad[13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[13]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N20
cycloneive_lcell_comb \temp_dMemLoad[12]~feeder (
// Equation(s):
// \temp_dMemLoad[12]~feeder_combout  = ramiframload_12

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_12),
	.cin(gnd),
	.combout(\temp_dMemLoad[12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[12]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N16
cycloneive_lcell_comb \temp_dMemLoad[10]~feeder (
// Equation(s):
// \temp_dMemLoad[10]~feeder_combout  = ramiframload_10

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_10),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_dMemLoad[10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[10]~feeder .lut_mask = 16'hF0F0;
defparam \temp_dMemLoad[10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N24
cycloneive_lcell_comb \temp_npc[10]~feeder (
// Equation(s):
// \temp_npc[10]~feeder_combout  = temp_npc_10

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_npc_101),
	.cin(gnd),
	.combout(\temp_npc[10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc[10]~feeder .lut_mask = 16'hFF00;
defparam \temp_npc[10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N30
cycloneive_lcell_comb \temp_dMemLoad[11]~feeder (
// Equation(s):
// \temp_dMemLoad[11]~feeder_combout  = ramiframload_11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_11),
	.cin(gnd),
	.combout(\temp_dMemLoad[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[11]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N10
cycloneive_lcell_comb \temp_dMemLoad[9]~feeder (
// Equation(s):
// \temp_dMemLoad[9]~feeder_combout  = ramiframload_9

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_9),
	.cin(gnd),
	.combout(\temp_dMemLoad[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[9]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N16
cycloneive_lcell_comb \temp_upper16[31]~feeder (
// Equation(s):
// \temp_upper16[31]~feeder_combout  = temp_iMemLoad_15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_iMemLoad_15),
	.cin(gnd),
	.combout(\temp_upper16[31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_upper16[31]~feeder .lut_mask = 16'hFF00;
defparam \temp_upper16[31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N20
cycloneive_lcell_comb \temp_dMemLoad[31]~feeder (
// Equation(s):
// \temp_dMemLoad[31]~feeder_combout  = ramiframload_31

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_31),
	.cin(gnd),
	.combout(\temp_dMemLoad[31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[31]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N12
cycloneive_lcell_comb \temp_dMemLoad[30]~feeder (
// Equation(s):
// \temp_dMemLoad[30]~feeder_combout  = ramiframload_30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_30),
	.cin(gnd),
	.combout(\temp_dMemLoad[30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[30]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N0
cycloneive_lcell_comb \temp_upper16[30]~feeder (
// Equation(s):
// \temp_upper16[30]~feeder_combout  = temp_iMemLoad_14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_iMemLoad_14),
	.cin(gnd),
	.combout(\temp_upper16[30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_upper16[30]~feeder .lut_mask = 16'hFF00;
defparam \temp_upper16[30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N6
cycloneive_lcell_comb \temp_upper16[29]~feeder (
// Equation(s):
// \temp_upper16[29]~feeder_combout  = temp_iMemLoad_13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_iMemLoad_13),
	.cin(gnd),
	.combout(\temp_upper16[29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_upper16[29]~feeder .lut_mask = 16'hFF00;
defparam \temp_upper16[29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N4
cycloneive_lcell_comb \temp_dMemLoad[29]~feeder (
// Equation(s):
// \temp_dMemLoad[29]~feeder_combout  = ramiframload_29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_29),
	.cin(gnd),
	.combout(\temp_dMemLoad[29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[29]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N8
cycloneive_lcell_comb \temp_dMemLoad[26]~feeder (
// Equation(s):
// \temp_dMemLoad[26]~feeder_combout  = ramiframload_26

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_26),
	.cin(gnd),
	.combout(\temp_dMemLoad[26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[26]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N16
cycloneive_lcell_comb \temp_dMemLoad[25]~feeder (
// Equation(s):
// \temp_dMemLoad[25]~feeder_combout  = ramiframload_25

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_dMemLoad[25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[25]~feeder .lut_mask = 16'hF0F0;
defparam \temp_dMemLoad[25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N30
cycloneive_lcell_comb \temp_upper16[25]~feeder (
// Equation(s):
// \temp_upper16[25]~feeder_combout  = temp_iMemLoad_9

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_iMemLoad_9),
	.cin(gnd),
	.combout(\temp_upper16[25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_upper16[25]~feeder .lut_mask = 16'hFF00;
defparam \temp_upper16[25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N8
cycloneive_lcell_comb \temp_npc[25]~feeder (
// Equation(s):
// \temp_npc[25]~feeder_combout  = temp_npc_25

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_npc_251),
	.cin(gnd),
	.combout(\temp_npc[25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc[25]~feeder .lut_mask = 16'hFF00;
defparam \temp_npc[25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N10
cycloneive_lcell_comb \temp_upper16[28]~feeder (
// Equation(s):
// \temp_upper16[28]~feeder_combout  = temp_iMemLoad_12

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_iMemLoad_12),
	.cin(gnd),
	.combout(\temp_upper16[28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_upper16[28]~feeder .lut_mask = 16'hFF00;
defparam \temp_upper16[28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N24
cycloneive_lcell_comb \temp_dMemLoad[27]~feeder (
// Equation(s):
// \temp_dMemLoad[27]~feeder_combout  = ramiframload_27

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_27),
	.cin(gnd),
	.combout(\temp_dMemLoad[27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[27]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N12
cycloneive_lcell_comb \temp_dMemLoad[17]~feeder (
// Equation(s):
// \temp_dMemLoad[17]~feeder_combout  = ramiframload_17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_17),
	.cin(gnd),
	.combout(\temp_dMemLoad[17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[17]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N24
cycloneive_lcell_comb \temp_npc[17]~feeder (
// Equation(s):
// \temp_npc[17]~feeder_combout  = temp_npc_17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_npc_171),
	.cin(gnd),
	.combout(\temp_npc[17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc[17]~feeder .lut_mask = 16'hFF00;
defparam \temp_npc[17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N10
cycloneive_lcell_comb \temp_dMemLoad[20]~feeder (
// Equation(s):
// \temp_dMemLoad[20]~feeder_combout  = ramiframload_20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_20),
	.cin(gnd),
	.combout(\temp_dMemLoad[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[20]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N2
cycloneive_lcell_comb \temp_npc[20]~feeder (
// Equation(s):
// \temp_npc[20]~feeder_combout  = temp_npc_20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_npc_201),
	.cin(gnd),
	.combout(\temp_npc[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc[20]~feeder .lut_mask = 16'hFF00;
defparam \temp_npc[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N24
cycloneive_lcell_comb \temp_upper16[19]~feeder (
// Equation(s):
// \temp_upper16[19]~feeder_combout  = temp_iMemLoad_3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_iMemLoad_3),
	.cin(gnd),
	.combout(\temp_upper16[19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_upper16[19]~feeder .lut_mask = 16'hFF00;
defparam \temp_upper16[19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N0
cycloneive_lcell_comb \temp_npc[19]~feeder (
// Equation(s):
// \temp_npc[19]~feeder_combout  = temp_npc_19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_npc_191),
	.cin(gnd),
	.combout(\temp_npc[19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_npc[19]~feeder .lut_mask = 16'hFF00;
defparam \temp_npc[19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N28
cycloneive_lcell_comb \temp_dMemLoad[18]~feeder (
// Equation(s):
// \temp_dMemLoad[18]~feeder_combout  = ramiframload_18

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_18),
	.datad(gnd),
	.cin(gnd),
	.combout(\temp_dMemLoad[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[18]~feeder .lut_mask = 16'hF0F0;
defparam \temp_dMemLoad[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N18
cycloneive_lcell_comb \temp_dMemLoad[24]~feeder (
// Equation(s):
// \temp_dMemLoad[24]~feeder_combout  = ramiframload_24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_24),
	.cin(gnd),
	.combout(\temp_dMemLoad[24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[24]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N16
cycloneive_lcell_comb \temp_dMemLoad[23]~feeder (
// Equation(s):
// \temp_dMemLoad[23]~feeder_combout  = ramiframload_23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_23),
	.cin(gnd),
	.combout(\temp_dMemLoad[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[23]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N12
cycloneive_lcell_comb \temp_upper16[23]~feeder (
// Equation(s):
// \temp_upper16[23]~feeder_combout  = temp_iMemLoad_7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_iMemLoad_7),
	.cin(gnd),
	.combout(\temp_upper16[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_upper16[23]~feeder .lut_mask = 16'hFF00;
defparam \temp_upper16[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N14
cycloneive_lcell_comb \temp_upper16[22]~feeder (
// Equation(s):
// \temp_upper16[22]~feeder_combout  = temp_iMemLoad_6

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_iMemLoad_6),
	.cin(gnd),
	.combout(\temp_upper16[22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_upper16[22]~feeder .lut_mask = 16'hFF00;
defparam \temp_upper16[22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N18
cycloneive_lcell_comb \temp_dMemLoad[22]~feeder (
// Equation(s):
// \temp_dMemLoad[22]~feeder_combout  = ramiframload_22

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_22),
	.cin(gnd),
	.combout(\temp_dMemLoad[22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[22]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N14
cycloneive_lcell_comb \temp_dMemLoad[21]~feeder (
// Equation(s):
// \temp_dMemLoad[21]~feeder_combout  = ramiframload_21

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_21),
	.cin(gnd),
	.combout(\temp_dMemLoad[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \temp_dMemLoad[21]~feeder .lut_mask = 16'hFF00;
defparam \temp_dMemLoad[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module npc_mux (
	temp_zeroFlag,
	branch_count_output_2,
	pc_count_four_output_2,
	pc_count_four_output_3,
	branch_count_output_3,
	pc_count_four_output_4,
	pc_count_four_output_5,
	branch_count_output_4,
	branch_count_output_5,
	pc_count_four_output_6,
	pc_count_four_output_7,
	branch_count_output_6,
	branch_count_output_7,
	pc_count_four_output_8,
	pc_count_four_output_9,
	branch_count_output_8,
	branch_count_output_9,
	pc_count_four_output_10,
	pc_count_four_output_11,
	branch_count_output_10,
	branch_count_output_11,
	pc_count_four_output_12,
	pc_count_four_output_13,
	branch_count_output_12,
	branch_count_output_13,
	pc_count_four_output_14,
	pc_count_four_output_15,
	branch_count_output_14,
	branch_count_output_15,
	pc_count_four_output_16,
	pc_count_four_output_17,
	branch_count_output_16,
	branch_count_output_17,
	pc_count_four_output_18,
	pc_count_four_output_19,
	branch_count_output_18,
	branch_count_output_19,
	branch_count_output_20,
	pc_count_four_output_20,
	pc_count_four_output_21,
	branch_count_output_21,
	pc_count_four_output_22,
	pc_count_four_output_23,
	branch_count_output_22,
	branch_count_output_23,
	pc_count_four_output_24,
	pc_count_four_output_25,
	branch_count_output_24,
	branch_count_output_25,
	branch_count_output_26,
	pc_count_four_output_26,
	pc_count_four_output_27,
	pc_count_four_output_28,
	branch_count_output_27,
	pc_count_four_output_29,
	branch_count_output_28,
	branch_count_output_29,
	pc_count_four_output_30,
	pc_count_four_output_31,
	branch_count_output_30,
	branch_count_output_31,
	pccount_1,
	pccount_0,
	temp_iMemLoad_0,
	temp_iMemLoad_15,
	temp_iMemLoad_14,
	temp_iMemLoad_13,
	temp_iMemLoad_10,
	temp_iMemLoad_9,
	temp_iMemLoad_12,
	temp_iMemLoad_11,
	temp_iMemLoad_1,
	temp_iMemLoad_4,
	temp_iMemLoad_3,
	temp_iMemLoad_2,
	temp_iMemLoad_8,
	temp_iMemLoad_7,
	temp_iMemLoad_6,
	temp_iMemLoad_5,
	temp_branchSelect,
	temp_rdat1_1,
	temp_npc_1,
	temp_pcselect_1,
	temp_pcselect_0,
	Mux30,
	temp_rdat1_0,
	temp_npc_0,
	Mux31,
	temp_rdat1_2,
	Mux29,
	temp_rdat1_3,
	Mux28,
	temp_rdat1_5,
	Mux26,
	temp_rdat1_4,
	Mux27,
	temp_rdat1_7,
	Mux24,
	temp_rdat1_6,
	Mux25,
	temp_rdat1_9,
	Mux22,
	temp_rdat1_8,
	Mux23,
	temp_rdat1_11,
	Mux20,
	temp_rdat1_10,
	Mux21,
	temp_rdat1_13,
	Mux18,
	temp_rdat1_12,
	Mux19,
	temp_rdat1_15,
	Mux16,
	temp_rdat1_14,
	Mux17,
	temp_rdat1_17,
	Mux14,
	temp_rdat1_16,
	Mux15,
	temp_rdat1_19,
	temp_iMemLoad_17,
	Mux12,
	temp_rdat1_18,
	temp_iMemLoad_16,
	Mux13,
	temp_rdat1_20,
	temp_iMemLoad_18,
	Mux11,
	temp_rdat1_21,
	temp_iMemLoad_19,
	Mux10,
	temp_rdat1_23,
	temp_iMemLoad_21,
	Mux8,
	temp_rdat1_22,
	temp_iMemLoad_20,
	Mux9,
	temp_rdat1_25,
	temp_iMemLoad_23,
	Mux6,
	temp_rdat1_24,
	temp_iMemLoad_22,
	Mux7,
	temp_rdat1_26,
	Mux5,
	temp_rdat1_27,
	Mux4,
	temp_rdat1_29,
	Mux2,
	temp_rdat1_28,
	Mux3,
	temp_rdat1_31,
	Mux0,
	temp_rdat1_30,
	Mux1,
	devpor,
	devclrn,
	devoe);
input 	temp_zeroFlag;
input 	branch_count_output_2;
input 	pc_count_four_output_2;
input 	pc_count_four_output_3;
input 	branch_count_output_3;
input 	pc_count_four_output_4;
input 	pc_count_four_output_5;
input 	branch_count_output_4;
input 	branch_count_output_5;
input 	pc_count_four_output_6;
input 	pc_count_four_output_7;
input 	branch_count_output_6;
input 	branch_count_output_7;
input 	pc_count_four_output_8;
input 	pc_count_four_output_9;
input 	branch_count_output_8;
input 	branch_count_output_9;
input 	pc_count_four_output_10;
input 	pc_count_four_output_11;
input 	branch_count_output_10;
input 	branch_count_output_11;
input 	pc_count_four_output_12;
input 	pc_count_four_output_13;
input 	branch_count_output_12;
input 	branch_count_output_13;
input 	pc_count_four_output_14;
input 	pc_count_four_output_15;
input 	branch_count_output_14;
input 	branch_count_output_15;
input 	pc_count_four_output_16;
input 	pc_count_four_output_17;
input 	branch_count_output_16;
input 	branch_count_output_17;
input 	pc_count_four_output_18;
input 	pc_count_four_output_19;
input 	branch_count_output_18;
input 	branch_count_output_19;
input 	branch_count_output_20;
input 	pc_count_four_output_20;
input 	pc_count_four_output_21;
input 	branch_count_output_21;
input 	pc_count_four_output_22;
input 	pc_count_four_output_23;
input 	branch_count_output_22;
input 	branch_count_output_23;
input 	pc_count_four_output_24;
input 	pc_count_four_output_25;
input 	branch_count_output_24;
input 	branch_count_output_25;
input 	branch_count_output_26;
input 	pc_count_four_output_26;
input 	pc_count_four_output_27;
input 	pc_count_four_output_28;
input 	branch_count_output_27;
input 	pc_count_four_output_29;
input 	branch_count_output_28;
input 	branch_count_output_29;
input 	pc_count_four_output_30;
input 	pc_count_four_output_31;
input 	branch_count_output_30;
input 	branch_count_output_31;
input 	pccount_1;
input 	pccount_0;
input 	temp_iMemLoad_0;
input 	temp_iMemLoad_15;
input 	temp_iMemLoad_14;
input 	temp_iMemLoad_13;
input 	temp_iMemLoad_10;
input 	temp_iMemLoad_9;
input 	temp_iMemLoad_12;
input 	temp_iMemLoad_11;
input 	temp_iMemLoad_1;
input 	temp_iMemLoad_4;
input 	temp_iMemLoad_3;
input 	temp_iMemLoad_2;
input 	temp_iMemLoad_8;
input 	temp_iMemLoad_7;
input 	temp_iMemLoad_6;
input 	temp_iMemLoad_5;
input 	temp_branchSelect;
input 	temp_rdat1_1;
input 	temp_npc_1;
input 	temp_pcselect_1;
input 	temp_pcselect_0;
output 	Mux30;
input 	temp_rdat1_0;
input 	temp_npc_0;
output 	Mux31;
input 	temp_rdat1_2;
output 	Mux29;
input 	temp_rdat1_3;
output 	Mux28;
input 	temp_rdat1_5;
output 	Mux26;
input 	temp_rdat1_4;
output 	Mux27;
input 	temp_rdat1_7;
output 	Mux24;
input 	temp_rdat1_6;
output 	Mux25;
input 	temp_rdat1_9;
output 	Mux22;
input 	temp_rdat1_8;
output 	Mux23;
input 	temp_rdat1_11;
output 	Mux20;
input 	temp_rdat1_10;
output 	Mux21;
input 	temp_rdat1_13;
output 	Mux18;
input 	temp_rdat1_12;
output 	Mux19;
input 	temp_rdat1_15;
output 	Mux16;
input 	temp_rdat1_14;
output 	Mux17;
input 	temp_rdat1_17;
output 	Mux14;
input 	temp_rdat1_16;
output 	Mux15;
input 	temp_rdat1_19;
input 	temp_iMemLoad_17;
output 	Mux12;
input 	temp_rdat1_18;
input 	temp_iMemLoad_16;
output 	Mux13;
input 	temp_rdat1_20;
input 	temp_iMemLoad_18;
output 	Mux11;
input 	temp_rdat1_21;
input 	temp_iMemLoad_19;
output 	Mux10;
input 	temp_rdat1_23;
input 	temp_iMemLoad_21;
output 	Mux8;
input 	temp_rdat1_22;
input 	temp_iMemLoad_20;
output 	Mux9;
input 	temp_rdat1_25;
input 	temp_iMemLoad_23;
output 	Mux6;
input 	temp_rdat1_24;
input 	temp_iMemLoad_22;
output 	Mux7;
input 	temp_rdat1_26;
output 	Mux5;
input 	temp_rdat1_27;
output 	Mux4;
input 	temp_rdat1_29;
output 	Mux2;
input 	temp_rdat1_28;
output 	Mux3;
input 	temp_rdat1_31;
output 	Mux0;
input 	temp_rdat1_30;
output 	Mux1;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Mux30~0_combout ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux29~0_combout ;
wire \Mux28~0_combout ;
wire \Mux26~0_combout ;
wire \Mux27~0_combout ;
wire \Mux24~0_combout ;
wire \Mux25~0_combout ;
wire \Mux22~0_combout ;
wire \Mux23~0_combout ;
wire \Mux20~0_combout ;
wire \Mux21~0_combout ;
wire \Mux18~0_combout ;
wire \Mux19~0_combout ;
wire \Mux16~0_combout ;
wire \Mux17~0_combout ;
wire \Mux14~0_combout ;
wire \Mux15~0_combout ;
wire \Mux12~0_combout ;
wire \Mux13~0_combout ;
wire \Mux11~0_combout ;
wire \Mux10~0_combout ;
wire \Mux8~0_combout ;
wire \Mux9~0_combout ;
wire \Mux6~0_combout ;
wire \Mux7~0_combout ;
wire \Mux5~0_combout ;
wire \Mux4~0_combout ;
wire \Mux2~0_combout ;
wire \Mux3~2_combout ;
wire \Mux0~0_combout ;
wire \Mux1~0_combout ;


// Location: LCCOMB_X62_Y42_N22
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// Mux30 = (\Mux31~0_combout  & ((pccount_1))) # (!\Mux31~0_combout  & (\Mux30~0_combout ))

	.dataa(\Mux30~0_combout ),
	.datab(pccount_1),
	.datac(gnd),
	.datad(\Mux31~0_combout ),
	.cin(gnd),
	.combout(Mux30),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hCCAA;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N18
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// Mux31 = (\Mux31~0_combout  & (pccount_0)) # (!\Mux31~0_combout  & ((\Mux31~1_combout )))

	.dataa(pccount_0),
	.datab(\Mux31~1_combout ),
	.datac(gnd),
	.datad(\Mux31~0_combout ),
	.cin(gnd),
	.combout(Mux31),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hAACC;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N20
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// Mux29 = (\Mux29~0_combout  & ((temp_iMemLoad_0) # ((!\Mux3~0_combout )))) # (!\Mux29~0_combout  & (((\branch_count_output[2]~0_combout  & \Mux3~0_combout ))))

	.dataa(\Mux29~0_combout ),
	.datab(temp_iMemLoad_0),
	.datac(branch_count_output_2),
	.datad(\Mux3~0_combout ),
	.cin(gnd),
	.combout(Mux29),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hD8AA;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N10
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// Mux28 = (\Mux28~0_combout  & (((temp_iMemLoad_1) # (!\Mux3~1_combout )))) # (!\Mux28~0_combout  & (\pc_count_four_output[3]~2_combout  & ((\Mux3~1_combout ))))

	.dataa(\Mux28~0_combout ),
	.datab(pc_count_four_output_3),
	.datac(temp_iMemLoad_1),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(Mux28),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hE4AA;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N8
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// Mux26 = (\Mux26~0_combout  & (((temp_iMemLoad_3) # (!\Mux3~1_combout )))) # (!\Mux26~0_combout  & (\pc_count_four_output[5]~6_combout  & ((\Mux3~1_combout ))))

	.dataa(\Mux26~0_combout ),
	.datab(pc_count_four_output_5),
	.datac(temp_iMemLoad_3),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(Mux26),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hE4AA;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N14
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// Mux27 = (\Mux3~0_combout  & ((\Mux27~0_combout  & (temp_iMemLoad_2)) # (!\Mux27~0_combout  & ((\branch_count_output[4]~4_combout ))))) # (!\Mux3~0_combout  & (((\Mux27~0_combout ))))

	.dataa(temp_iMemLoad_2),
	.datab(\Mux3~0_combout ),
	.datac(branch_count_output_4),
	.datad(\Mux27~0_combout ),
	.cin(gnd),
	.combout(Mux27),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hBBC0;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N16
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// Mux24 = (\Mux24~0_combout  & (((temp_iMemLoad_5)) # (!\Mux3~1_combout ))) # (!\Mux24~0_combout  & (\Mux3~1_combout  & ((\pc_count_four_output[7]~10_combout ))))

	.dataa(\Mux24~0_combout ),
	.datab(\Mux3~1_combout ),
	.datac(temp_iMemLoad_5),
	.datad(pc_count_four_output_7),
	.cin(gnd),
	.combout(Mux24),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hE6A2;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y45_N0
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// Mux25 = (\Mux25~0_combout  & ((temp_iMemLoad_4) # ((!\Mux3~0_combout )))) # (!\Mux25~0_combout  & (((\Mux3~0_combout  & \branch_count_output[6]~8_combout ))))

	.dataa(\Mux25~0_combout ),
	.datab(temp_iMemLoad_4),
	.datac(\Mux3~0_combout ),
	.datad(branch_count_output_6),
	.cin(gnd),
	.combout(Mux25),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hDA8A;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N30
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// Mux22 = (\Mux3~1_combout  & ((\Mux22~0_combout  & ((temp_iMemLoad_7))) # (!\Mux22~0_combout  & (\pc_count_four_output[9]~14_combout )))) # (!\Mux3~1_combout  & (((\Mux22~0_combout ))))

	.dataa(pc_count_four_output_9),
	.datab(temp_iMemLoad_7),
	.datac(\Mux3~1_combout ),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(Mux22),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hCFA0;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N18
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// Mux23 = (\Mux3~0_combout  & ((\Mux23~0_combout  & ((temp_iMemLoad_6))) # (!\Mux23~0_combout  & (\branch_count_output[8]~12_combout )))) # (!\Mux3~0_combout  & (((\Mux23~0_combout ))))

	.dataa(branch_count_output_8),
	.datab(\Mux3~0_combout ),
	.datac(temp_iMemLoad_6),
	.datad(\Mux23~0_combout ),
	.cin(gnd),
	.combout(Mux23),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hF388;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N20
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// Mux20 = (\Mux20~0_combout  & ((temp_iMemLoad_9) # ((!\Mux3~1_combout )))) # (!\Mux20~0_combout  & (((\pc_count_four_output[11]~18_combout  & \Mux3~1_combout ))))

	.dataa(\Mux20~0_combout ),
	.datab(temp_iMemLoad_9),
	.datac(pc_count_four_output_11),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(Mux20),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hD8AA;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N20
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// Mux21 = (\Mux21~0_combout  & ((temp_iMemLoad_8) # ((!\Mux3~1_combout )))) # (!\Mux21~0_combout  & (((\pc_count_four_output[10]~16_combout  & \Mux3~1_combout ))))

	.dataa(temp_iMemLoad_8),
	.datab(pc_count_four_output_10),
	.datac(\Mux21~0_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(Mux21),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hACF0;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N8
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// Mux18 = (\Mux18~0_combout  & ((temp_iMemLoad_11) # ((!\Mux3~1_combout )))) # (!\Mux18~0_combout  & (((\pc_count_four_output[13]~22_combout  & \Mux3~1_combout ))))

	.dataa(temp_iMemLoad_11),
	.datab(pc_count_four_output_13),
	.datac(\Mux18~0_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(Mux18),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hACF0;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N30
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// Mux19 = (\Mux3~0_combout  & ((\Mux19~0_combout  & (temp_iMemLoad_10)) # (!\Mux19~0_combout  & ((\branch_count_output[12]~20_combout ))))) # (!\Mux3~0_combout  & (((\Mux19~0_combout ))))

	.dataa(temp_iMemLoad_10),
	.datab(branch_count_output_12),
	.datac(\Mux3~0_combout ),
	.datad(\Mux19~0_combout ),
	.cin(gnd),
	.combout(Mux19),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hAFC0;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N14
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// Mux16 = (\Mux16~0_combout  & (((temp_iMemLoad_13) # (!\Mux3~1_combout )))) # (!\Mux16~0_combout  & (\pc_count_four_output[15]~26_combout  & ((\Mux3~1_combout ))))

	.dataa(pc_count_four_output_15),
	.datab(\Mux16~0_combout ),
	.datac(temp_iMemLoad_13),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(Mux16),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hE2CC;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N30
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// Mux17 = (\Mux17~0_combout  & (((temp_iMemLoad_12)) # (!\Mux3~0_combout ))) # (!\Mux17~0_combout  & (\Mux3~0_combout  & ((\branch_count_output[14]~24_combout ))))

	.dataa(\Mux17~0_combout ),
	.datab(\Mux3~0_combout ),
	.datac(temp_iMemLoad_12),
	.datad(branch_count_output_14),
	.cin(gnd),
	.combout(Mux17),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hE6A2;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N12
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// Mux14 = (\Mux14~0_combout  & (((temp_iMemLoad_15) # (!\Mux3~1_combout )))) # (!\Mux14~0_combout  & (\pc_count_four_output[17]~30_combout  & ((\Mux3~1_combout ))))

	.dataa(\Mux14~0_combout ),
	.datab(pc_count_four_output_17),
	.datac(temp_iMemLoad_15),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(Mux14),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hE4AA;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y46_N8
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// Mux15 = (\Mux3~0_combout  & ((\Mux15~0_combout  & ((temp_iMemLoad_14))) # (!\Mux15~0_combout  & (\branch_count_output[16]~28_combout )))) # (!\Mux3~0_combout  & (((\Mux15~0_combout ))))

	.dataa(branch_count_output_16),
	.datab(\Mux3~0_combout ),
	.datac(temp_iMemLoad_14),
	.datad(\Mux15~0_combout ),
	.cin(gnd),
	.combout(Mux15),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hF388;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y46_N12
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// Mux12 = (\Mux3~1_combout  & ((\Mux12~0_combout  & (temp_iMemLoad_17)) # (!\Mux12~0_combout  & ((\pc_count_four_output[19]~34_combout ))))) # (!\Mux3~1_combout  & (((\Mux12~0_combout ))))

	.dataa(\Mux3~1_combout ),
	.datab(temp_iMemLoad_17),
	.datac(pc_count_four_output_19),
	.datad(\Mux12~0_combout ),
	.cin(gnd),
	.combout(Mux12),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hDDA0;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y40_N18
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// Mux13 = (\Mux3~0_combout  & ((\Mux13~0_combout  & ((temp_iMemLoad_16))) # (!\Mux13~0_combout  & (\branch_count_output[18]~32_combout )))) # (!\Mux3~0_combout  & (((\Mux13~0_combout ))))

	.dataa(\Mux3~0_combout ),
	.datab(branch_count_output_18),
	.datac(temp_iMemLoad_16),
	.datad(\Mux13~0_combout ),
	.cin(gnd),
	.combout(Mux13),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hF588;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N4
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// Mux11 = (\Mux11~0_combout  & (((temp_iMemLoad_18)) # (!\Mux3~0_combout ))) # (!\Mux11~0_combout  & (\Mux3~0_combout  & (\branch_count_output[20]~36_combout )))

	.dataa(\Mux11~0_combout ),
	.datab(\Mux3~0_combout ),
	.datac(branch_count_output_20),
	.datad(temp_iMemLoad_18),
	.cin(gnd),
	.combout(Mux11),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hEA62;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N2
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// Mux10 = (\Mux3~1_combout  & ((\Mux10~0_combout  & (temp_iMemLoad_19)) # (!\Mux10~0_combout  & ((\pc_count_four_output[21]~38_combout ))))) # (!\Mux3~1_combout  & (((\Mux10~0_combout ))))

	.dataa(\Mux3~1_combout ),
	.datab(temp_iMemLoad_19),
	.datac(\Mux10~0_combout ),
	.datad(pc_count_four_output_21),
	.cin(gnd),
	.combout(Mux10),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hDAD0;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N24
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// Mux8 = (\Mux3~1_combout  & ((\Mux8~0_combout  & ((temp_iMemLoad_21))) # (!\Mux8~0_combout  & (\pc_count_four_output[23]~42_combout )))) # (!\Mux3~1_combout  & (((\Mux8~0_combout ))))

	.dataa(\Mux3~1_combout ),
	.datab(pc_count_four_output_23),
	.datac(temp_iMemLoad_21),
	.datad(\Mux8~0_combout ),
	.cin(gnd),
	.combout(Mux8),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hF588;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N4
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// Mux9 = (\Mux9~0_combout  & (((temp_iMemLoad_20) # (!\Mux3~0_combout )))) # (!\Mux9~0_combout  & (\branch_count_output[22]~40_combout  & (\Mux3~0_combout )))

	.dataa(branch_count_output_22),
	.datab(\Mux9~0_combout ),
	.datac(\Mux3~0_combout ),
	.datad(temp_iMemLoad_20),
	.cin(gnd),
	.combout(Mux9),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hEC2C;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N12
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// Mux6 = (\Mux3~1_combout  & ((\Mux6~0_combout  & (temp_iMemLoad_23)) # (!\Mux6~0_combout  & ((\pc_count_four_output[25]~46_combout ))))) # (!\Mux3~1_combout  & (\Mux6~0_combout ))

	.dataa(\Mux3~1_combout ),
	.datab(\Mux6~0_combout ),
	.datac(temp_iMemLoad_23),
	.datad(pc_count_four_output_25),
	.cin(gnd),
	.combout(Mux6),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hE6C4;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N28
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// Mux7 = (\Mux3~0_combout  & ((\Mux7~0_combout  & (temp_iMemLoad_22)) # (!\Mux7~0_combout  & ((\branch_count_output[24]~44_combout ))))) # (!\Mux3~0_combout  & (((\Mux7~0_combout ))))

	.dataa(temp_iMemLoad_22),
	.datab(\Mux3~0_combout ),
	.datac(branch_count_output_24),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(Mux7),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hBBC0;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N24
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// Mux5 = (\Mux5~0_combout  & ((\pc_count_four_output[28]~52_combout ) # ((!\Mux3~0_combout )))) # (!\Mux5~0_combout  & (((\Mux3~0_combout  & \branch_count_output[26]~48_combout ))))

	.dataa(\Mux5~0_combout ),
	.datab(pc_count_four_output_28),
	.datac(\Mux3~0_combout ),
	.datad(branch_count_output_26),
	.cin(gnd),
	.combout(Mux5),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hDA8A;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y46_N14
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// Mux4 = (\Mux3~0_combout  & ((\Mux4~0_combout  & ((\pc_count_four_output[29]~54_combout ))) # (!\Mux4~0_combout  & (\branch_count_output[27]~50_combout )))) # (!\Mux3~0_combout  & (((\Mux4~0_combout ))))

	.dataa(branch_count_output_27),
	.datab(pc_count_four_output_29),
	.datac(\Mux3~0_combout ),
	.datad(\Mux4~0_combout ),
	.cin(gnd),
	.combout(Mux4),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hCFA0;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y46_N26
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// Mux2 = (\Mux3~1_combout  & ((\Mux2~0_combout  & ((\pc_count_four_output[31]~58_combout ))) # (!\Mux2~0_combout  & (\pc_count_four_output[29]~54_combout )))) # (!\Mux3~1_combout  & (((\Mux2~0_combout ))))

	.dataa(\Mux3~1_combout ),
	.datab(pc_count_four_output_29),
	.datac(\Mux2~0_combout ),
	.datad(pc_count_four_output_31),
	.cin(gnd),
	.combout(Mux2),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hF858;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N28
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// Mux3 = (\Mux3~2_combout  & ((\pc_count_four_output[30]~56_combout ) # ((!\Mux3~0_combout )))) # (!\Mux3~2_combout  & (((\Mux3~0_combout  & \branch_count_output[28]~52_combout ))))

	.dataa(\Mux3~2_combout ),
	.datab(pc_count_four_output_30),
	.datac(\Mux3~0_combout ),
	.datad(branch_count_output_28),
	.cin(gnd),
	.combout(Mux3),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hDA8A;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N14
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// Mux0 = (\Mux31~0_combout  & (\pc_count_four_output[31]~58_combout )) # (!\Mux31~0_combout  & ((\Mux0~0_combout )))

	.dataa(gnd),
	.datab(\Mux31~0_combout ),
	.datac(pc_count_four_output_31),
	.datad(\Mux0~0_combout ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hF3C0;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N8
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// Mux1 = (\Mux31~0_combout  & (\pc_count_four_output[30]~56_combout )) # (!\Mux31~0_combout  & ((\Mux1~0_combout )))

	.dataa(gnd),
	.datab(\Mux31~0_combout ),
	.datac(pc_count_four_output_30),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(Mux1),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hF3C0;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N10
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (temp_pcselect_1 & (((!temp_pcselect_0 & temp_npc_1)))) # (!temp_pcselect_1 & (temp_rdat1_1))

	.dataa(temp_rdat1_1),
	.datab(temp_pcselect_0),
	.datac(temp_pcselect_1),
	.datad(temp_npc_1),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'h3A0A;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N20
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (!temp_pcselect_0 & ((temp_zeroFlag1 $ (temp_branchSelect1)) # (!temp_pcselect_1)))

	.dataa(temp_zeroFlag),
	.datab(temp_branchSelect),
	.datac(temp_pcselect_1),
	.datad(temp_pcselect_0),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'h006F;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N0
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (temp_pcselect_1 & (!temp_pcselect_0 & ((temp_npc_0)))) # (!temp_pcselect_1 & (((temp_rdat1_0))))

	.dataa(temp_pcselect_1),
	.datab(temp_pcselect_0),
	.datac(temp_rdat1_0),
	.datad(temp_npc_0),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'h7250;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N4
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (temp_pcselect_1 & ((temp_pcselect_0) # (temp_zeroFlag1 $ (!temp_branchSelect1))))

	.dataa(temp_zeroFlag),
	.datab(temp_branchSelect),
	.datac(temp_pcselect_1),
	.datad(temp_pcselect_0),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hF090;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N6
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (temp_pcselect_1 & ((temp_pcselect_0) # (temp_zeroFlag1 $ (temp_branchSelect1)))) # (!temp_pcselect_1 & (((!temp_pcselect_0))))

	.dataa(temp_zeroFlag),
	.datab(temp_branchSelect),
	.datac(temp_pcselect_1),
	.datad(temp_pcselect_0),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hF06F;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N6
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (\Mux3~0_combout  & (((\Mux3~1_combout )))) # (!\Mux3~0_combout  & ((\Mux3~1_combout  & ((\pc_count_four_output[2]~0_combout ))) # (!\Mux3~1_combout  & (temp_rdat1_2))))

	.dataa(\Mux3~0_combout ),
	.datab(temp_rdat1_2),
	.datac(pc_count_four_output_2),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hFA44;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N12
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (\Mux3~0_combout  & ((\branch_count_output[3]~2_combout ) # ((\Mux3~1_combout )))) # (!\Mux3~0_combout  & (((temp_rdat1_3 & !\Mux3~1_combout ))))

	.dataa(\Mux3~0_combout ),
	.datab(branch_count_output_3),
	.datac(temp_rdat1_3),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hAAD8;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N6
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (\Mux3~1_combout  & (((\Mux3~0_combout )))) # (!\Mux3~1_combout  & ((\Mux3~0_combout  & (\branch_count_output[5]~6_combout )) # (!\Mux3~0_combout  & ((temp_rdat1_5)))))

	.dataa(\Mux3~1_combout ),
	.datab(branch_count_output_5),
	.datac(\Mux3~0_combout ),
	.datad(temp_rdat1_5),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hE5E0;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y44_N12
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (\Mux3~0_combout  & (((\Mux3~1_combout )))) # (!\Mux3~0_combout  & ((\Mux3~1_combout  & ((\pc_count_four_output[4]~4_combout ))) # (!\Mux3~1_combout  & (temp_rdat1_4))))

	.dataa(temp_rdat1_4),
	.datab(\Mux3~0_combout ),
	.datac(\Mux3~1_combout ),
	.datad(pc_count_four_output_4),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hF2C2;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N6
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (\Mux3~0_combout  & ((\Mux3~1_combout ) # ((\branch_count_output[7]~10_combout )))) # (!\Mux3~0_combout  & (!\Mux3~1_combout  & ((temp_rdat1_7))))

	.dataa(\Mux3~0_combout ),
	.datab(\Mux3~1_combout ),
	.datac(branch_count_output_7),
	.datad(temp_rdat1_7),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hB9A8;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N28
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (\Mux3~0_combout  & (((\Mux3~1_combout )))) # (!\Mux3~0_combout  & ((\Mux3~1_combout  & (\pc_count_four_output[6]~8_combout )) # (!\Mux3~1_combout  & ((temp_rdat1_6)))))

	.dataa(pc_count_four_output_6),
	.datab(temp_rdat1_6),
	.datac(\Mux3~0_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hFA0C;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N20
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (\Mux3~1_combout  & (((\Mux3~0_combout )))) # (!\Mux3~1_combout  & ((\Mux3~0_combout  & ((\branch_count_output[9]~14_combout ))) # (!\Mux3~0_combout  & (temp_rdat1_9))))

	.dataa(temp_rdat1_9),
	.datab(\Mux3~1_combout ),
	.datac(\Mux3~0_combout ),
	.datad(branch_count_output_9),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hF2C2;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N12
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (\Mux3~0_combout  & (((\Mux3~1_combout )))) # (!\Mux3~0_combout  & ((\Mux3~1_combout  & ((\pc_count_four_output[8]~12_combout ))) # (!\Mux3~1_combout  & (temp_rdat1_8))))

	.dataa(temp_rdat1_8),
	.datab(\Mux3~0_combout ),
	.datac(pc_count_four_output_8),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hFC22;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N10
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (\Mux3~1_combout  & (((\Mux3~0_combout )))) # (!\Mux3~1_combout  & ((\Mux3~0_combout  & ((\branch_count_output[11]~18_combout ))) # (!\Mux3~0_combout  & (temp_rdat1_11))))

	.dataa(\Mux3~1_combout ),
	.datab(temp_rdat1_11),
	.datac(\Mux3~0_combout ),
	.datad(branch_count_output_11),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hF4A4;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N14
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (\Mux3~0_combout  & ((\branch_count_output[10]~16_combout ) # ((\Mux3~1_combout )))) # (!\Mux3~0_combout  & (((temp_rdat1_10 & !\Mux3~1_combout ))))

	.dataa(branch_count_output_10),
	.datab(temp_rdat1_10),
	.datac(\Mux3~0_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hF0AC;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N22
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (\Mux3~1_combout  & (((\Mux3~0_combout )))) # (!\Mux3~1_combout  & ((\Mux3~0_combout  & ((\branch_count_output[13]~22_combout ))) # (!\Mux3~0_combout  & (temp_rdat1_13))))

	.dataa(\Mux3~1_combout ),
	.datab(temp_rdat1_13),
	.datac(\Mux3~0_combout ),
	.datad(branch_count_output_13),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hF4A4;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N24
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (\Mux3~1_combout  & (((\Mux3~0_combout ) # (\pc_count_four_output[12]~20_combout )))) # (!\Mux3~1_combout  & (temp_rdat1_12 & (!\Mux3~0_combout )))

	.dataa(\Mux3~1_combout ),
	.datab(temp_rdat1_12),
	.datac(\Mux3~0_combout ),
	.datad(pc_count_four_output_12),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hAEA4;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N0
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (\Mux3~0_combout  & ((\Mux3~1_combout ) # ((\branch_count_output[15]~26_combout )))) # (!\Mux3~0_combout  & (!\Mux3~1_combout  & ((temp_rdat1_15))))

	.dataa(\Mux3~0_combout ),
	.datab(\Mux3~1_combout ),
	.datac(branch_count_output_15),
	.datad(temp_rdat1_15),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hB9A8;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N12
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (\Mux3~0_combout  & (((\Mux3~1_combout )))) # (!\Mux3~0_combout  & ((\Mux3~1_combout  & (\pc_count_four_output[14]~24_combout )) # (!\Mux3~1_combout  & ((temp_rdat1_14)))))

	.dataa(pc_count_four_output_14),
	.datab(temp_rdat1_14),
	.datac(\Mux3~0_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hFA0C;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y46_N0
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (\Mux3~1_combout  & (((\Mux3~0_combout )))) # (!\Mux3~1_combout  & ((\Mux3~0_combout  & ((\branch_count_output[17]~30_combout ))) # (!\Mux3~0_combout  & (temp_rdat1_17))))

	.dataa(\Mux3~1_combout ),
	.datab(temp_rdat1_17),
	.datac(\Mux3~0_combout ),
	.datad(branch_count_output_17),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hF4A4;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y46_N2
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (\Mux3~1_combout  & ((\pc_count_four_output[16]~28_combout ) # ((\Mux3~0_combout )))) # (!\Mux3~1_combout  & (((!\Mux3~0_combout  & temp_rdat1_16))))

	.dataa(\Mux3~1_combout ),
	.datab(pc_count_four_output_16),
	.datac(\Mux3~0_combout ),
	.datad(temp_rdat1_16),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hADA8;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y46_N10
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (\Mux3~0_combout  & (((\branch_count_output[19]~34_combout ) # (\Mux3~1_combout )))) # (!\Mux3~0_combout  & (temp_rdat1_19 & ((!\Mux3~1_combout ))))

	.dataa(temp_rdat1_19),
	.datab(\Mux3~0_combout ),
	.datac(branch_count_output_19),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hCCE2;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N16
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (\Mux3~0_combout  & (((\Mux3~1_combout )))) # (!\Mux3~0_combout  & ((\Mux3~1_combout  & (\pc_count_four_output[18]~32_combout )) # (!\Mux3~1_combout  & ((temp_rdat1_18)))))

	.dataa(pc_count_four_output_18),
	.datab(\Mux3~0_combout ),
	.datac(temp_rdat1_18),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hEE30;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y45_N10
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (\Mux3~0_combout  & (((\Mux3~1_combout )))) # (!\Mux3~0_combout  & ((\Mux3~1_combout  & ((\pc_count_four_output[20]~36_combout ))) # (!\Mux3~1_combout  & (temp_rdat1_20))))

	.dataa(temp_rdat1_20),
	.datab(pc_count_four_output_20),
	.datac(\Mux3~0_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hFC0A;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N30
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (\Mux3~0_combout  & ((\branch_count_output[21]~38_combout ) # ((\Mux3~1_combout )))) # (!\Mux3~0_combout  & (((temp_rdat1_21 & !\Mux3~1_combout ))))

	.dataa(\Mux3~0_combout ),
	.datab(branch_count_output_21),
	.datac(temp_rdat1_21),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hAAD8;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N0
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (\Mux3~1_combout  & (\Mux3~0_combout )) # (!\Mux3~1_combout  & ((\Mux3~0_combout  & (\branch_count_output[23]~42_combout )) # (!\Mux3~0_combout  & ((temp_rdat1_23)))))

	.dataa(\Mux3~1_combout ),
	.datab(\Mux3~0_combout ),
	.datac(branch_count_output_23),
	.datad(temp_rdat1_23),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hD9C8;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N20
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (\Mux3~1_combout  & ((\pc_count_four_output[22]~40_combout ) # ((\Mux3~0_combout )))) # (!\Mux3~1_combout  & (((!\Mux3~0_combout  & temp_rdat1_22))))

	.dataa(pc_count_four_output_22),
	.datab(\Mux3~1_combout ),
	.datac(\Mux3~0_combout ),
	.datad(temp_rdat1_22),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hCBC8;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N10
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (\Mux3~0_combout  & ((\Mux3~1_combout ) # ((\branch_count_output[25]~46_combout )))) # (!\Mux3~0_combout  & (!\Mux3~1_combout  & (temp_rdat1_25)))

	.dataa(\Mux3~0_combout ),
	.datab(\Mux3~1_combout ),
	.datac(temp_rdat1_25),
	.datad(branch_count_output_25),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hBA98;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N16
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (\Mux3~1_combout  & (((\pc_count_four_output[24]~44_combout ) # (\Mux3~0_combout )))) # (!\Mux3~1_combout  & (temp_rdat1_24 & ((!\Mux3~0_combout ))))

	.dataa(\Mux3~1_combout ),
	.datab(temp_rdat1_24),
	.datac(pc_count_four_output_24),
	.datad(\Mux3~0_combout ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hAAE4;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N6
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (\Mux3~0_combout  & (((\Mux3~1_combout )))) # (!\Mux3~0_combout  & ((\Mux3~1_combout  & ((\pc_count_four_output[26]~48_combout ))) # (!\Mux3~1_combout  & (temp_rdat1_26))))

	.dataa(\Mux3~0_combout ),
	.datab(temp_rdat1_26),
	.datac(pc_count_four_output_26),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hFA44;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N16
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (\Mux3~0_combout  & (((\Mux3~1_combout )))) # (!\Mux3~0_combout  & ((\Mux3~1_combout  & (\pc_count_four_output[27]~50_combout )) # (!\Mux3~1_combout  & ((temp_rdat1_27)))))

	.dataa(pc_count_four_output_27),
	.datab(temp_rdat1_27),
	.datac(\Mux3~0_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hFA0C;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y46_N4
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (\Mux3~1_combout  & (\Mux3~0_combout )) # (!\Mux3~1_combout  & ((\Mux3~0_combout  & ((\branch_count_output[29]~54_combout ))) # (!\Mux3~0_combout  & (temp_rdat1_29))))

	.dataa(\Mux3~1_combout ),
	.datab(\Mux3~0_combout ),
	.datac(temp_rdat1_29),
	.datad(branch_count_output_29),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hDC98;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y44_N26
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (\Mux3~0_combout  & (((\Mux3~1_combout )))) # (!\Mux3~0_combout  & ((\Mux3~1_combout  & ((\pc_count_four_output[28]~52_combout ))) # (!\Mux3~1_combout  & (temp_rdat1_28))))

	.dataa(temp_rdat1_28),
	.datab(pc_count_four_output_28),
	.datac(\Mux3~0_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hFC0A;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N28
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (temp_pcselect_1 & (((\branch_count_output[31]~58_combout  & !temp_pcselect_0)))) # (!temp_pcselect_1 & (temp_rdat1_31))

	.dataa(temp_rdat1_31),
	.datab(branch_count_output_31),
	.datac(temp_pcselect_1),
	.datad(temp_pcselect_0),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'h0ACA;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N2
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (temp_pcselect_1 & (\branch_count_output[30]~56_combout  & (!temp_pcselect_0))) # (!temp_pcselect_1 & (((temp_rdat1_30))))

	.dataa(branch_count_output_30),
	.datab(temp_pcselect_0),
	.datac(temp_pcselect_1),
	.datad(temp_rdat1_30),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'h2F20;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module program_count (
	pccount_1,
	pccount_0,
	pccount_2,
	pccount_3,
	pccount_5,
	pccount_4,
	pccount_7,
	pccount_6,
	pccount_9,
	pccount_8,
	pccount_11,
	pccount_10,
	pccount_13,
	pccount_12,
	pccount_15,
	pccount_14,
	pccount_17,
	pccount_16,
	pccount_19,
	pccount_18,
	pccount_20,
	pccount_21,
	pccount_23,
	pccount_22,
	pccount_25,
	pccount_24,
	pccount_26,
	pccount_27,
	pccount_29,
	pccount_28,
	pccount_31,
	pccount_30,
	Mux30,
	wen,
	Mux31,
	Mux29,
	Mux28,
	Mux26,
	Mux27,
	Mux24,
	Mux25,
	Mux22,
	Mux23,
	Mux20,
	Mux21,
	Mux18,
	Mux19,
	Mux16,
	Mux17,
	Mux14,
	Mux15,
	Mux12,
	Mux13,
	Mux11,
	Mux10,
	Mux8,
	Mux9,
	Mux6,
	Mux7,
	Mux5,
	Mux4,
	Mux2,
	Mux3,
	Mux0,
	Mux1,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	pccount_1;
output 	pccount_0;
output 	pccount_2;
output 	pccount_3;
output 	pccount_5;
output 	pccount_4;
output 	pccount_7;
output 	pccount_6;
output 	pccount_9;
output 	pccount_8;
output 	pccount_11;
output 	pccount_10;
output 	pccount_13;
output 	pccount_12;
output 	pccount_15;
output 	pccount_14;
output 	pccount_17;
output 	pccount_16;
output 	pccount_19;
output 	pccount_18;
output 	pccount_20;
output 	pccount_21;
output 	pccount_23;
output 	pccount_22;
output 	pccount_25;
output 	pccount_24;
output 	pccount_26;
output 	pccount_27;
output 	pccount_29;
output 	pccount_28;
output 	pccount_31;
output 	pccount_30;
input 	Mux30;
input 	wen;
input 	Mux31;
input 	Mux29;
input 	Mux28;
input 	Mux26;
input 	Mux27;
input 	Mux24;
input 	Mux25;
input 	Mux22;
input 	Mux23;
input 	Mux20;
input 	Mux21;
input 	Mux18;
input 	Mux19;
input 	Mux16;
input 	Mux17;
input 	Mux14;
input 	Mux15;
input 	Mux12;
input 	Mux13;
input 	Mux11;
input 	Mux10;
input 	Mux8;
input 	Mux9;
input 	Mux6;
input 	Mux7;
input 	Mux5;
input 	Mux4;
input 	Mux2;
input 	Mux3;
input 	Mux0;
input 	Mux1;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: FF_X63_Y43_N13
dffeas \pccount[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_1),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[1] .is_wysiwyg = "true";
defparam \pccount[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y43_N29
dffeas \pccount[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_0),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[0] .is_wysiwyg = "true";
defparam \pccount[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N21
dffeas \pccount[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_2),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[2] .is_wysiwyg = "true";
defparam \pccount[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N13
dffeas \pccount[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_3),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[3] .is_wysiwyg = "true";
defparam \pccount[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N31
dffeas \pccount[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_5),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[5] .is_wysiwyg = "true";
defparam \pccount[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N9
dffeas \pccount[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_4),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[4] .is_wysiwyg = "true";
defparam \pccount[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N9
dffeas \pccount[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_7),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[7] .is_wysiwyg = "true";
defparam \pccount[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N11
dffeas \pccount[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_6),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[6] .is_wysiwyg = "true";
defparam \pccount[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N11
dffeas \pccount[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_9),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[9] .is_wysiwyg = "true";
defparam \pccount[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N1
dffeas \pccount[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_8),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[8] .is_wysiwyg = "true";
defparam \pccount[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y43_N1
dffeas \pccount[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_11),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[11] .is_wysiwyg = "true";
defparam \pccount[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y43_N7
dffeas \pccount[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_10),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[10] .is_wysiwyg = "true";
defparam \pccount[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y43_N15
dffeas \pccount[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_13),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[13] .is_wysiwyg = "true";
defparam \pccount[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y43_N3
dffeas \pccount[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_12),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[12] .is_wysiwyg = "true";
defparam \pccount[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N11
dffeas \pccount[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_15),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[15] .is_wysiwyg = "true";
defparam \pccount[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N17
dffeas \pccount[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_14),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[14] .is_wysiwyg = "true";
defparam \pccount[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y43_N27
dffeas \pccount[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_17),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[17] .is_wysiwyg = "true";
defparam \pccount[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y43_N19
dffeas \pccount[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_16),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[16] .is_wysiwyg = "true";
defparam \pccount[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y43_N3
dffeas \pccount[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_19),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[19] .is_wysiwyg = "true";
defparam \pccount[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y43_N13
dffeas \pccount[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_18),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[18] .is_wysiwyg = "true";
defparam \pccount[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y43_N19
dffeas \pccount[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_20),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[20] .is_wysiwyg = "true";
defparam \pccount[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N31
dffeas \pccount[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_21),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[21] .is_wysiwyg = "true";
defparam \pccount[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N5
dffeas \pccount[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_23),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[23] .is_wysiwyg = "true";
defparam \pccount[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N29
dffeas \pccount[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_22),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[22] .is_wysiwyg = "true";
defparam \pccount[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y43_N5
dffeas \pccount[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_25),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[25] .is_wysiwyg = "true";
defparam \pccount[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y43_N21
dffeas \pccount[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_24),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[24] .is_wysiwyg = "true";
defparam \pccount[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y43_N9
dffeas \pccount[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_26),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[26] .is_wysiwyg = "true";
defparam \pccount[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y43_N29
dffeas \pccount[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_27),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[27] .is_wysiwyg = "true";
defparam \pccount[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N1
dffeas \pccount[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_29),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[29] .is_wysiwyg = "true";
defparam \pccount[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y43_N1
dffeas \pccount[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_28),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[28] .is_wysiwyg = "true";
defparam \pccount[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N29
dffeas \pccount[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_31),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[31] .is_wysiwyg = "true";
defparam \pccount[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y43_N9
dffeas \pccount[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(wen),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pccount_30),
	.prn(vcc));
// synopsys translate_off
defparam \pccount[30] .is_wysiwyg = "true";
defparam \pccount[30] .power_up = "low";
// synopsys translate_on

endmodule

module register_file (
	temp_regwrite,
	temp_branchDest_1,
	temp_branchDest_0,
	temp_branchDest_3,
	temp_branchDest_2,
	temp_branchDest_4,
	Mux30,
	Mux31,
	Mux29,
	Mux27,
	Mux28,
	Mux23,
	Mux24,
	Mux25,
	Mux26,
	Mux15,
	Mux17,
	Mux16,
	Mux18,
	Mux19,
	Mux21,
	Mux20,
	Mux22,
	Mux0,
	Mux1,
	Mux2,
	Mux5,
	Mux6,
	Mux3,
	Mux4,
	Mux14,
	Mux11,
	Mux12,
	Mux13,
	Mux7,
	Mux8,
	Mux9,
	Mux10,
	temp_imemload_output_17,
	temp_imemload_output_16,
	temp_imemload_output_19,
	temp_imemload_output_18,
	temp_imemload_output_22,
	temp_imemload_output_21,
	temp_imemload_output_24,
	temp_imemload_output_23,
	Mux62,
	Mux621,
	Mux301,
	Mux302,
	Mux63,
	Mux631,
	Mux311,
	Mux312,
	Mux291,
	Mux292,
	Mux271,
	Mux272,
	Mux281,
	Mux282,
	Mux61,
	Mux611,
	Mux231,
	Mux232,
	Mux241,
	Mux242,
	Mux251,
	Mux252,
	Mux261,
	Mux262,
	Mux60,
	Mux601,
	Mux151,
	Mux152,
	Mux171,
	Mux172,
	Mux161,
	Mux162,
	Mux181,
	Mux182,
	Mux191,
	Mux192,
	Mux211,
	Mux212,
	Mux201,
	Mux202,
	Mux221,
	Mux222,
	Mux59,
	Mux591,
	Mux01,
	Mux02,
	Mux110,
	Mux111,
	Mux210,
	Mux213,
	Mux51,
	Mux52,
	Mux64,
	Mux65,
	Mux32,
	Mux33,
	Mux41,
	Mux42,
	Mux141,
	Mux142,
	Mux112,
	Mux113,
	Mux121,
	Mux122,
	Mux131,
	Mux132,
	Mux71,
	Mux72,
	Mux81,
	Mux82,
	Mux91,
	Mux92,
	Mux101,
	Mux102,
	Mux48,
	Mux481,
	Mux511,
	Mux512,
	Mux36,
	Mux361,
	Mux45,
	Mux451,
	Mux46,
	Mux461,
	Mux47,
	Mux471,
	Mux321,
	Mux322,
	Mux331,
	Mux332,
	Mux34,
	Mux341,
	Mux35,
	Mux351,
	Mux37,
	Mux371,
	Mux38,
	Mux381,
	Mux39,
	Mux391,
	Mux40,
	Mux401,
	Mux411,
	Mux412,
	Mux421,
	Mux422,
	Mux43,
	Mux431,
	Mux44,
	Mux441,
	Mux53,
	Mux531,
	Mux49,
	Mux491,
	Mux54,
	Mux541,
	Mux55,
	Mux551,
	Mux56,
	Mux561,
	Mux57,
	Mux571,
	Mux58,
	Mux581,
	Mux50,
	Mux501,
	Mux521,
	Mux522,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	temp_regwrite;
input 	temp_branchDest_1;
input 	temp_branchDest_0;
input 	temp_branchDest_3;
input 	temp_branchDest_2;
input 	temp_branchDest_4;
input 	Mux30;
input 	Mux31;
input 	Mux29;
input 	Mux27;
input 	Mux28;
input 	Mux23;
input 	Mux24;
input 	Mux25;
input 	Mux26;
input 	Mux15;
input 	Mux17;
input 	Mux16;
input 	Mux18;
input 	Mux19;
input 	Mux21;
input 	Mux20;
input 	Mux22;
input 	Mux0;
input 	Mux1;
input 	Mux2;
input 	Mux5;
input 	Mux6;
input 	Mux3;
input 	Mux4;
input 	Mux14;
input 	Mux11;
input 	Mux12;
input 	Mux13;
input 	Mux7;
input 	Mux8;
input 	Mux9;
input 	Mux10;
input 	temp_imemload_output_17;
input 	temp_imemload_output_16;
input 	temp_imemload_output_19;
input 	temp_imemload_output_18;
input 	temp_imemload_output_22;
input 	temp_imemload_output_21;
input 	temp_imemload_output_24;
input 	temp_imemload_output_23;
output 	Mux62;
output 	Mux621;
output 	Mux301;
output 	Mux302;
output 	Mux63;
output 	Mux631;
output 	Mux311;
output 	Mux312;
output 	Mux291;
output 	Mux292;
output 	Mux271;
output 	Mux272;
output 	Mux281;
output 	Mux282;
output 	Mux61;
output 	Mux611;
output 	Mux231;
output 	Mux232;
output 	Mux241;
output 	Mux242;
output 	Mux251;
output 	Mux252;
output 	Mux261;
output 	Mux262;
output 	Mux60;
output 	Mux601;
output 	Mux151;
output 	Mux152;
output 	Mux171;
output 	Mux172;
output 	Mux161;
output 	Mux162;
output 	Mux181;
output 	Mux182;
output 	Mux191;
output 	Mux192;
output 	Mux211;
output 	Mux212;
output 	Mux201;
output 	Mux202;
output 	Mux221;
output 	Mux222;
output 	Mux59;
output 	Mux591;
output 	Mux01;
output 	Mux02;
output 	Mux110;
output 	Mux111;
output 	Mux210;
output 	Mux213;
output 	Mux51;
output 	Mux52;
output 	Mux64;
output 	Mux65;
output 	Mux32;
output 	Mux33;
output 	Mux41;
output 	Mux42;
output 	Mux141;
output 	Mux142;
output 	Mux112;
output 	Mux113;
output 	Mux121;
output 	Mux122;
output 	Mux131;
output 	Mux132;
output 	Mux71;
output 	Mux72;
output 	Mux81;
output 	Mux82;
output 	Mux91;
output 	Mux92;
output 	Mux101;
output 	Mux102;
output 	Mux48;
output 	Mux481;
output 	Mux511;
output 	Mux512;
output 	Mux36;
output 	Mux361;
output 	Mux45;
output 	Mux451;
output 	Mux46;
output 	Mux461;
output 	Mux47;
output 	Mux471;
output 	Mux321;
output 	Mux322;
output 	Mux331;
output 	Mux332;
output 	Mux34;
output 	Mux341;
output 	Mux35;
output 	Mux351;
output 	Mux37;
output 	Mux371;
output 	Mux38;
output 	Mux381;
output 	Mux39;
output 	Mux391;
output 	Mux40;
output 	Mux401;
output 	Mux411;
output 	Mux412;
output 	Mux421;
output 	Mux422;
output 	Mux43;
output 	Mux431;
output 	Mux44;
output 	Mux441;
output 	Mux53;
output 	Mux531;
output 	Mux49;
output 	Mux491;
output 	Mux54;
output 	Mux541;
output 	Mux55;
output 	Mux551;
output 	Mux56;
output 	Mux561;
output 	Mux57;
output 	Mux571;
output 	Mux58;
output 	Mux581;
output 	Mux50;
output 	Mux501;
output 	Mux521;
output 	Mux522;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \storeregister[22][1]~q ;
wire \storeregister[18][1]~q ;
wire \Mux62~2_combout ;
wire \Mux62~12_combout ;
wire \Mux30~2_combout ;
wire \Mux30~4_combout ;
wire \Mux30~14_combout ;
wire \storeregister[26][0]~q ;
wire \storeregister[18][0]~q ;
wire \Mux63~2_combout ;
wire \Mux63~4_combout ;
wire \Mux63~12_combout ;
wire \storeregister[1][0]~q ;
wire \Mux63~14_combout ;
wire \Mux31~2_combout ;
wire \storeregister[28][2]~q ;
wire \storeregister[30][3]~q ;
wire \Mux28~14_combout ;
wire \storeregister[16][8]~q ;
wire \Mux23~4_combout ;
wire \Mux23~12_combout ;
wire \Mux23~14_combout ;
wire \storeregister[26][7]~q ;
wire \Mux25~12_combout ;
wire \storeregister[8][5]~q ;
wire \Mux26~12_combout ;
wire \Mux17~12_combout ;
wire \Mux17~14_combout ;
wire \Mux16~4_combout ;
wire \Mux16~12_combout ;
wire \storeregister[20][13]~q ;
wire \Mux18~4_combout ;
wire \storeregister[8][13]~q ;
wire \Mux18~12_combout ;
wire \Mux19~12_combout ;
wire \Mux21~4_combout ;
wire \storeregister[30][11]~q ;
wire \storeregister[8][11]~q ;
wire \Mux20~12_combout ;
wire \storeregister[1][11]~q ;
wire \storeregister[18][9]~q ;
wire \Mux22~2_combout ;
wire \Mux22~4_combout ;
wire \Mux59~2_combout ;
wire \Mux59~4_combout ;
wire \Mux59~12_combout ;
wire \storeregister[18][31]~q ;
wire \Mux0~2_combout ;
wire \storeregister[8][31]~q ;
wire \Mux0~12_combout ;
wire \storeregister[1][31]~q ;
wire \storeregister[4][30]~q ;
wire \Mux1~12_combout ;
wire \Mux2~14_combout ;
wire \Mux5~12_combout ;
wire \storeregister[26][25]~q ;
wire \storeregister[4][25]~q ;
wire \storeregister[8][25]~q ;
wire \Mux6~12_combout ;
wire \storeregister[28][28]~q ;
wire \storeregister[8][28]~q ;
wire \storeregister[4][28]~q ;
wire \Mux3~12_combout ;
wire \Mux4~2_combout ;
wire \storeregister[18][17]~q ;
wire \Mux14~2_combout ;
wire \storeregister[20][17]~q ;
wire \storeregister[16][20]~q ;
wire \Mux11~4_combout ;
wire \Mux11~14_combout ;
wire \storeregister[8][19]~q ;
wire \Mux12~12_combout ;
wire \storeregister[18][18]~q ;
wire \Mux13~2_combout ;
wire \storeregister[3][18]~q ;
wire \storeregister[1][18]~q ;
wire \Mux13~14_combout ;
wire \storeregister[22][24]~q ;
wire \Mux8~2_combout ;
wire \Mux8~12_combout ;
wire \storeregister[26][22]~q ;
wire \storeregister[18][22]~q ;
wire \Mux9~2_combout ;
wire \Mux9~14_combout ;
wire \Mux10~4_combout ;
wire \Mux48~2_combout ;
wire \Mux36~14_combout ;
wire \Mux45~2_combout ;
wire \Mux45~14_combout ;
wire \Mux46~2_combout ;
wire \Mux47~4_combout ;
wire \Mux32~2_combout ;
wire \Mux32~14_combout ;
wire \Mux34~2_combout ;
wire \Mux34~4_combout ;
wire \Mux34~12_combout ;
wire \Mux35~12_combout ;
wire \Mux38~2_combout ;
wire \Mux38~12_combout ;
wire \Mux39~2_combout ;
wire \Mux40~12_combout ;
wire \Mux42~2_combout ;
wire \Mux43~2_combout ;
wire \Mux49~4_combout ;
wire \Mux54~2_combout ;
wire \Mux55~4_combout ;
wire \Mux56~2_combout ;
wire \Mux56~12_combout ;
wire \Mux57~4_combout ;
wire \Mux58~2_combout ;
wire \Mux50~2_combout ;
wire \Mux52~14_combout ;
wire \Decoder0~13_combout ;
wire \Decoder0~20_combout ;
wire \storeregister[18][1]~feeder_combout ;
wire \storeregister[28][2]~feeder_combout ;
wire \storeregister[30][3]~feeder_combout ;
wire \storeregister[20][13]~feeder_combout ;
wire \storeregister[30][11]~feeder_combout ;
wire \storeregister[18][31]~feeder_combout ;
wire \storeregister[26][25]~feeder_combout ;
wire \storeregister[28][28]~feeder_combout ;
wire \storeregister[20][17]~feeder_combout ;
wire \storeregister[22][24]~feeder_combout ;
wire \storeregister[26][22]~feeder_combout ;
wire \storeregister[31][1]~feeder_combout ;
wire \Decoder0~9_combout ;
wire \Decoder0~27_combout ;
wire \storeregister[31][1]~q ;
wire \storeregister[27][1]~feeder_combout ;
wire \Decoder0~25_combout ;
wire \storeregister[27][1]~q ;
wire \storeregister[19][1]~feeder_combout ;
wire \Decoder0~26_combout ;
wire \storeregister[19][1]~q ;
wire \Mux62~7_combout ;
wire \storeregister[23][1]~feeder_combout ;
wire \Decoder0~24_combout ;
wire \storeregister[23][1]~q ;
wire \Mux62~8_combout ;
wire \storeregister[17][1]~feeder_combout ;
wire \Decoder0~44_combout ;
wire \storeregister[17][1]~q ;
wire \storeregister[25][1]~feeder_combout ;
wire \Decoder0~10_combout ;
wire \Decoder0~11_combout ;
wire \storeregister[25][1]~q ;
wire \Mux62~0_combout ;
wire \Decoder0~43_combout ;
wire \storeregister[21][1]~q ;
wire \storeregister[29][1]~feeder_combout ;
wire \Decoder0~12_combout ;
wire \storeregister[29][1]~q ;
wire \Mux62~1_combout ;
wire \storeregister[26][1]~feeder_combout ;
wire \Decoder0~14_combout ;
wire \storeregister[26][1]~q ;
wire \storeregister[30][1]~feeder_combout ;
wire \Decoder0~17_combout ;
wire \storeregister[30][1]~q ;
wire \Mux62~3_combout ;
wire \Decoder0~8_combout ;
wire \Decoder0~21_combout ;
wire \storeregister[20][1]~q ;
wire \Decoder0~22_combout ;
wire \storeregister[16][1]~q ;
wire \Mux62~4_combout ;
wire \storeregister[24][1]~feeder_combout ;
wire \Decoder0~19_combout ;
wire \storeregister[24][1]~q ;
wire \Mux62~5_combout ;
wire \Mux62~6_combout ;
wire \Decoder0~30_combout ;
wire \Decoder0~45_combout ;
wire \storeregister[5][1]~q ;
wire \Mux62~10_combout ;
wire \storeregister[7][1]~feeder_combout ;
wire \Decoder0~32_combout ;
wire \storeregister[7][1]~q ;
wire \storeregister[6][1]~feeder_combout ;
wire \Decoder0~28_combout ;
wire \Decoder0~29_combout ;
wire \storeregister[6][1]~q ;
wire \Mux62~11_combout ;
wire \Decoder0~42_combout ;
wire \storeregister[15][1]~q ;
wire \Decoder0~39_combout ;
wire \storeregister[14][1]~q ;
wire \Decoder0~40_combout ;
wire \storeregister[13][1]~q ;
wire \Decoder0~41_combout ;
wire \storeregister[12][1]~q ;
wire \Mux62~17_combout ;
wire \Mux62~18_combout ;
wire \storeregister[2][1]~feeder_combout ;
wire \Decoder0~38_combout ;
wire \storeregister[2][1]~q ;
wire \Decoder0~46_combout ;
wire \storeregister[1][1]~q ;
wire \Decoder0~37_combout ;
wire \storeregister[3][1]~q ;
wire \Mux62~14_combout ;
wire \Mux62~15_combout ;
wire \storeregister[11][1]~feeder_combout ;
wire \Decoder0~36_combout ;
wire \storeregister[11][1]~q ;
wire \Decoder0~33_combout ;
wire \storeregister[9][1]~q ;
wire \Mux62~13_combout ;
wire \Mux62~16_combout ;
wire \storeregister[28][1]~feeder_combout ;
wire \Decoder0~23_combout ;
wire \storeregister[28][1]~q ;
wire \Mux30~5_combout ;
wire \Mux30~3_combout ;
wire \Mux30~6_combout ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \Mux30~7_combout ;
wire \Mux30~8_combout ;
wire \Decoder0~31_combout ;
wire \storeregister[4][1]~q ;
wire \Mux30~10_combout ;
wire \Mux30~11_combout ;
wire \Decoder0~34_combout ;
wire \storeregister[10][1]~q ;
wire \storeregister[8][1]~feeder_combout ;
wire \Decoder0~18_combout ;
wire \Decoder0~35_combout ;
wire \storeregister[8][1]~q ;
wire \Mux30~12_combout ;
wire \Mux30~13_combout ;
wire \Mux30~15_combout ;
wire \Mux30~16_combout ;
wire \Mux30~17_combout ;
wire \Mux30~18_combout ;
wire \storeregister[29][0]~feeder_combout ;
wire \storeregister[29][0]~q ;
wire \storeregister[25][0]~feeder_combout ;
wire \storeregister[25][0]~q ;
wire \storeregister[21][0]~q ;
wire \storeregister[17][0]~q ;
wire \Mux63~0_combout ;
wire \Mux63~1_combout ;
wire \storeregister[30][0]~q ;
wire \Decoder0~15_combout ;
wire \storeregister[22][0]~q ;
wire \Mux63~3_combout ;
wire \storeregister[20][0]~q ;
wire \storeregister[28][0]~q ;
wire \Mux63~5_combout ;
wire \Mux63~6_combout ;
wire \storeregister[23][0]~feeder_combout ;
wire \storeregister[23][0]~q ;
wire \Mux63~7_combout ;
wire \storeregister[27][0]~feeder_combout ;
wire \storeregister[27][0]~q ;
wire \storeregister[31][0]~feeder_combout ;
wire \storeregister[31][0]~q ;
wire \Mux63~8_combout ;
wire \storeregister[10][0]~q ;
wire \Mux63~10_combout ;
wire \storeregister[11][0]~q ;
wire \storeregister[9][0]~q ;
wire \Mux63~11_combout ;
wire \storeregister[6][0]~feeder_combout ;
wire \storeregister[6][0]~q ;
wire \storeregister[7][0]~feeder_combout ;
wire \storeregister[7][0]~q ;
wire \Mux63~13_combout ;
wire \storeregister[2][0]~q ;
wire \Mux63~15_combout ;
wire \Mux63~16_combout ;
wire \storeregister[15][0]~feeder_combout ;
wire \storeregister[15][0]~q ;
wire \storeregister[12][0]~feeder_combout ;
wire \storeregister[12][0]~q ;
wire \storeregister[13][0]~feeder_combout ;
wire \storeregister[13][0]~q ;
wire \Mux63~17_combout ;
wire \storeregister[14][0]~feeder_combout ;
wire \storeregister[14][0]~q ;
wire \Mux63~18_combout ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \storeregister[19][0]~feeder_combout ;
wire \storeregister[19][0]~q ;
wire \Mux31~7_combout ;
wire \Mux31~8_combout ;
wire \storeregister[24][0]~q ;
wire \storeregister[16][0]~q ;
wire \Mux31~4_combout ;
wire \Mux31~5_combout ;
wire \Mux31~3_combout ;
wire \Mux31~6_combout ;
wire \storeregister[3][0]~q ;
wire \Mux31~14_combout ;
wire \Mux31~15_combout ;
wire \storeregister[5][0]~q ;
wire \storeregister[4][0]~q ;
wire \Mux31~12_combout ;
wire \Mux31~13_combout ;
wire \Mux31~16_combout ;
wire \storeregister[8][0]~feeder_combout ;
wire \storeregister[8][0]~q ;
wire \Mux31~10_combout ;
wire \Mux31~11_combout ;
wire \Mux31~17_combout ;
wire \Mux31~18_combout ;
wire \storeregister[20][2]~q ;
wire \storeregister[16][2]~q ;
wire \storeregister[24][2]~feeder_combout ;
wire \storeregister[24][2]~q ;
wire \Mux29~4_combout ;
wire \Mux29~5_combout ;
wire \storeregister[30][2]~feeder_combout ;
wire \storeregister[30][2]~q ;
wire \storeregister[18][2]~feeder_combout ;
wire \Decoder0~16_combout ;
wire \storeregister[18][2]~q ;
wire \storeregister[26][2]~q ;
wire \Mux29~2_combout ;
wire \Mux29~3_combout ;
wire \Mux29~6_combout ;
wire \storeregister[19][2]~q ;
wire \storeregister[23][2]~q ;
wire \Mux29~7_combout ;
wire \storeregister[31][2]~feeder_combout ;
wire \storeregister[31][2]~q ;
wire \storeregister[27][2]~feeder_combout ;
wire \storeregister[27][2]~q ;
wire \Mux29~8_combout ;
wire \storeregister[25][2]~q ;
wire \storeregister[29][2]~q ;
wire \storeregister[17][2]~q ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \storeregister[5][2]~q ;
wire \storeregister[4][2]~q ;
wire \Mux29~12_combout ;
wire \storeregister[6][2]~feeder_combout ;
wire \storeregister[6][2]~q ;
wire \Mux29~13_combout ;
wire \storeregister[3][2]~q ;
wire \storeregister[1][2]~q ;
wire \Mux29~14_combout ;
wire \Mux29~15_combout ;
wire \Mux29~16_combout ;
wire \storeregister[12][2]~q ;
wire \storeregister[13][2]~q ;
wire \Mux29~17_combout ;
wire \storeregister[14][2]~feeder_combout ;
wire \storeregister[14][2]~q ;
wire \storeregister[15][2]~feeder_combout ;
wire \storeregister[15][2]~q ;
wire \Mux29~18_combout ;
wire \storeregister[9][2]~q ;
wire \storeregister[10][2]~q ;
wire \storeregister[8][2]~feeder_combout ;
wire \storeregister[8][2]~q ;
wire \Mux29~10_combout ;
wire \storeregister[11][2]~q ;
wire \Mux29~11_combout ;
wire \storeregister[31][4]~feeder_combout ;
wire \storeregister[31][4]~q ;
wire \storeregister[27][4]~q ;
wire \storeregister[23][4]~q ;
wire \storeregister[19][4]~q ;
wire \Mux27~7_combout ;
wire \Mux27~8_combout ;
wire \storeregister[16][4]~q ;
wire \storeregister[24][4]~feeder_combout ;
wire \storeregister[24][4]~q ;
wire \Mux27~4_combout ;
wire \storeregister[20][4]~q ;
wire \storeregister[28][4]~q ;
wire \Mux27~5_combout ;
wire \storeregister[26][4]~q ;
wire \storeregister[18][4]~feeder_combout ;
wire \storeregister[18][4]~q ;
wire \Mux27~2_combout ;
wire \storeregister[22][4]~q ;
wire \storeregister[30][4]~feeder_combout ;
wire \storeregister[30][4]~q ;
wire \Mux27~3_combout ;
wire \Mux27~6_combout ;
wire \storeregister[17][4]~q ;
wire \storeregister[21][4]~q ;
wire \Mux27~0_combout ;
wire \storeregister[29][4]~q ;
wire \storeregister[25][4]~q ;
wire \Mux27~1_combout ;
wire \storeregister[3][4]~q ;
wire \storeregister[1][4]~q ;
wire \Mux27~14_combout ;
wire \Mux27~15_combout ;
wire \storeregister[7][4]~feeder_combout ;
wire \storeregister[7][4]~q ;
wire \storeregister[4][4]~q ;
wire \storeregister[5][4]~q ;
wire \Mux27~12_combout ;
wire \Mux27~13_combout ;
wire \Mux27~16_combout ;
wire \storeregister[10][4]~q ;
wire \storeregister[8][4]~feeder_combout ;
wire \storeregister[8][4]~q ;
wire \Mux27~10_combout ;
wire \storeregister[9][4]~q ;
wire \storeregister[11][4]~feeder_combout ;
wire \storeregister[11][4]~q ;
wire \Mux27~11_combout ;
wire \storeregister[12][4]~q ;
wire \storeregister[13][4]~q ;
wire \Mux27~17_combout ;
wire \storeregister[14][4]~feeder_combout ;
wire \storeregister[14][4]~q ;
wire \storeregister[15][4]~feeder_combout ;
wire \storeregister[15][4]~q ;
wire \Mux27~18_combout ;
wire \storeregister[20][3]~q ;
wire \storeregister[16][3]~q ;
wire \Mux28~4_combout ;
wire \storeregister[28][3]~feeder_combout ;
wire \storeregister[28][3]~q ;
wire \Mux28~5_combout ;
wire \storeregister[22][3]~feeder_combout ;
wire \storeregister[22][3]~q ;
wire \storeregister[18][3]~q ;
wire \Mux28~2_combout ;
wire \storeregister[26][3]~q ;
wire \Mux28~3_combout ;
wire \Mux28~6_combout ;
wire \storeregister[25][3]~feeder_combout ;
wire \storeregister[25][3]~q ;
wire \storeregister[17][3]~q ;
wire \Mux28~0_combout ;
wire \storeregister[29][3]~q ;
wire \storeregister[21][3]~q ;
wire \Mux28~1_combout ;
wire \storeregister[27][3]~feeder_combout ;
wire \storeregister[27][3]~q ;
wire \Mux28~7_combout ;
wire \storeregister[23][3]~q ;
wire \storeregister[31][3]~feeder_combout ;
wire \storeregister[31][3]~q ;
wire \Mux28~8_combout ;
wire \storeregister[6][3]~feeder_combout ;
wire \storeregister[6][3]~q ;
wire \storeregister[5][3]~q ;
wire \storeregister[4][3]~q ;
wire \Mux28~10_combout ;
wire \storeregister[7][3]~feeder_combout ;
wire \storeregister[7][3]~q ;
wire \Mux28~11_combout ;
wire \storeregister[9][3]~feeder_combout ;
wire \storeregister[9][3]~q ;
wire \storeregister[11][3]~q ;
wire \storeregister[10][3]~q ;
wire \storeregister[8][3]~q ;
wire \Mux28~12_combout ;
wire \Mux28~13_combout ;
wire \storeregister[2][3]~q ;
wire \Mux28~15_combout ;
wire \Mux28~16_combout ;
wire \storeregister[15][3]~q ;
wire \storeregister[14][3]~q ;
wire \storeregister[12][3]~q ;
wire \storeregister[13][3]~q ;
wire \Mux28~17_combout ;
wire \Mux28~18_combout ;
wire \Mux61~4_combout ;
wire \Mux61~5_combout ;
wire \storeregister[22][2]~q ;
wire \Mux61~2_combout ;
wire \Mux61~3_combout ;
wire \Mux61~6_combout ;
wire \storeregister[21][2]~q ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \Mux61~7_combout ;
wire \Mux61~8_combout ;
wire \Mux61~14_combout ;
wire \storeregister[2][2]~feeder_combout ;
wire \storeregister[2][2]~q ;
wire \Mux61~15_combout ;
wire \Mux61~12_combout ;
wire \Mux61~13_combout ;
wire \Mux61~16_combout ;
wire \storeregister[7][2]~feeder_combout ;
wire \storeregister[7][2]~q ;
wire \Mux61~10_combout ;
wire \Mux61~11_combout ;
wire \Mux61~17_combout ;
wire \Mux61~18_combout ;
wire \storeregister[23][8]~q ;
wire \storeregister[19][8]~q ;
wire \Mux23~7_combout ;
wire \storeregister[27][8]~feeder_combout ;
wire \storeregister[27][8]~q ;
wire \storeregister[31][8]~feeder_combout ;
wire \storeregister[31][8]~q ;
wire \Mux23~8_combout ;
wire \storeregister[26][8]~q ;
wire \storeregister[18][8]~feeder_combout ;
wire \storeregister[18][8]~q ;
wire \Mux23~2_combout ;
wire \storeregister[30][8]~feeder_combout ;
wire \storeregister[30][8]~q ;
wire \Mux23~3_combout ;
wire \storeregister[28][8]~feeder_combout ;
wire \storeregister[28][8]~q ;
wire \storeregister[20][8]~feeder_combout ;
wire \storeregister[20][8]~q ;
wire \Mux23~5_combout ;
wire \Mux23~6_combout ;
wire \storeregister[21][8]~feeder_combout ;
wire \storeregister[21][8]~q ;
wire \storeregister[17][8]~feeder_combout ;
wire \storeregister[17][8]~q ;
wire \Mux23~0_combout ;
wire \storeregister[25][8]~q ;
wire \storeregister[29][8]~feeder_combout ;
wire \storeregister[29][8]~q ;
wire \Mux23~1_combout ;
wire \storeregister[11][8]~q ;
wire \storeregister[9][8]~q ;
wire \storeregister[8][8]~q ;
wire \storeregister[10][8]~q ;
wire \Mux23~10_combout ;
wire \Mux23~11_combout ;
wire \storeregister[7][8]~q ;
wire \storeregister[6][8]~q ;
wire \Mux23~13_combout ;
wire \storeregister[2][8]~q ;
wire \Mux23~15_combout ;
wire \Mux23~16_combout ;
wire \storeregister[14][8]~feeder_combout ;
wire \storeregister[14][8]~q ;
wire \storeregister[12][8]~q ;
wire \storeregister[13][8]~q ;
wire \Mux23~17_combout ;
wire \storeregister[15][8]~q ;
wire \Mux23~18_combout ;
wire \storeregister[25][7]~q ;
wire \storeregister[17][7]~feeder_combout ;
wire \storeregister[17][7]~q ;
wire \Mux24~0_combout ;
wire \storeregister[29][7]~feeder_combout ;
wire \storeregister[29][7]~q ;
wire \storeregister[21][7]~feeder_combout ;
wire \storeregister[21][7]~q ;
wire \Mux24~1_combout ;
wire \storeregister[23][7]~feeder_combout ;
wire \storeregister[23][7]~q ;
wire \storeregister[27][7]~feeder_combout ;
wire \storeregister[27][7]~q ;
wire \storeregister[19][7]~q ;
wire \Mux24~7_combout ;
wire \storeregister[31][7]~feeder_combout ;
wire \storeregister[31][7]~q ;
wire \Mux24~8_combout ;
wire \storeregister[22][7]~q ;
wire \storeregister[18][7]~q ;
wire \Mux24~2_combout ;
wire \storeregister[30][7]~feeder_combout ;
wire \storeregister[30][7]~q ;
wire \Mux24~3_combout ;
wire \storeregister[24][7]~feeder_combout ;
wire \storeregister[24][7]~q ;
wire \storeregister[28][7]~q ;
wire \storeregister[16][7]~q ;
wire \storeregister[20][7]~feeder_combout ;
wire \storeregister[20][7]~q ;
wire \Mux24~4_combout ;
wire \Mux24~5_combout ;
wire \Mux24~6_combout ;
wire \storeregister[6][7]~q ;
wire \storeregister[5][7]~q ;
wire \storeregister[4][7]~q ;
wire \Mux24~10_combout ;
wire \storeregister[7][7]~feeder_combout ;
wire \storeregister[7][7]~q ;
wire \Mux24~11_combout ;
wire \storeregister[14][7]~feeder_combout ;
wire \storeregister[14][7]~q ;
wire \storeregister[15][7]~q ;
wire \storeregister[13][7]~q ;
wire \storeregister[12][7]~q ;
wire \Mux24~17_combout ;
wire \Mux24~18_combout ;
wire \storeregister[8][7]~q ;
wire \storeregister[10][7]~q ;
wire \Mux24~12_combout ;
wire \storeregister[9][7]~feeder_combout ;
wire \storeregister[9][7]~q ;
wire \Mux24~13_combout ;
wire \storeregister[3][7]~q ;
wire \storeregister[1][7]~q ;
wire \Mux24~14_combout ;
wire \storeregister[2][7]~q ;
wire \Mux24~15_combout ;
wire \Mux24~16_combout ;
wire \storeregister[28][6]~feeder_combout ;
wire \storeregister[28][6]~q ;
wire \storeregister[16][6]~feeder_combout ;
wire \storeregister[16][6]~q ;
wire \storeregister[24][6]~feeder_combout ;
wire \storeregister[24][6]~q ;
wire \Mux25~4_combout ;
wire \storeregister[20][6]~feeder_combout ;
wire \storeregister[20][6]~q ;
wire \Mux25~5_combout ;
wire \storeregister[22][6]~q ;
wire \storeregister[30][6]~q ;
wire \storeregister[26][6]~q ;
wire \storeregister[18][6]~q ;
wire \Mux25~2_combout ;
wire \Mux25~3_combout ;
wire \Mux25~6_combout ;
wire \storeregister[23][6]~feeder_combout ;
wire \storeregister[23][6]~q ;
wire \storeregister[19][6]~feeder_combout ;
wire \storeregister[19][6]~q ;
wire \Mux25~7_combout ;
wire \storeregister[27][6]~feeder_combout ;
wire \storeregister[27][6]~q ;
wire \storeregister[31][6]~feeder_combout ;
wire \storeregister[31][6]~q ;
wire \Mux25~8_combout ;
wire \storeregister[21][6]~q ;
wire \Mux25~0_combout ;
wire \storeregister[25][6]~q ;
wire \storeregister[29][6]~feeder_combout ;
wire \storeregister[29][6]~q ;
wire \Mux25~1_combout ;
wire \storeregister[11][6]~q ;
wire \storeregister[10][6]~q ;
wire \storeregister[8][6]~q ;
wire \Mux25~10_combout ;
wire \storeregister[9][6]~q ;
wire \Mux25~11_combout ;
wire \storeregister[7][6]~q ;
wire \storeregister[6][6]~q ;
wire \Mux25~13_combout ;
wire \storeregister[3][6]~q ;
wire \storeregister[1][6]~q ;
wire \Mux25~14_combout ;
wire \storeregister[2][6]~feeder_combout ;
wire \storeregister[2][6]~q ;
wire \Mux25~15_combout ;
wire \Mux25~16_combout ;
wire \storeregister[15][6]~feeder_combout ;
wire \storeregister[15][6]~q ;
wire \storeregister[13][6]~q ;
wire \storeregister[12][6]~q ;
wire \Mux25~17_combout ;
wire \storeregister[14][6]~feeder_combout ;
wire \storeregister[14][6]~q ;
wire \Mux25~18_combout ;
wire \storeregister[18][5]~feeder_combout ;
wire \storeregister[18][5]~q ;
wire \Mux26~2_combout ;
wire \storeregister[26][5]~feeder_combout ;
wire \storeregister[26][5]~q ;
wire \Mux26~3_combout ;
wire \storeregister[28][5]~q ;
wire \storeregister[20][5]~feeder_combout ;
wire \storeregister[20][5]~q ;
wire \Mux26~4_combout ;
wire \Mux26~5_combout ;
wire \Mux26~6_combout ;
wire \storeregister[31][5]~q ;
wire \storeregister[23][5]~q ;
wire \storeregister[19][5]~q ;
wire \storeregister[27][5]~q ;
wire \Mux26~7_combout ;
wire \Mux26~8_combout ;
wire \storeregister[17][5]~feeder_combout ;
wire \storeregister[17][5]~q ;
wire \storeregister[25][5]~feeder_combout ;
wire \storeregister[25][5]~q ;
wire \Mux26~0_combout ;
wire \storeregister[21][5]~feeder_combout ;
wire \storeregister[21][5]~q ;
wire \storeregister[29][5]~feeder_combout ;
wire \storeregister[29][5]~q ;
wire \Mux26~1_combout ;
wire \storeregister[11][5]~q ;
wire \storeregister[9][5]~q ;
wire \Mux26~13_combout ;
wire \storeregister[2][5]~q ;
wire \storeregister[1][5]~q ;
wire \storeregister[3][5]~q ;
wire \Mux26~14_combout ;
wire \Mux26~15_combout ;
wire \Mux26~16_combout ;
wire \storeregister[14][5]~feeder_combout ;
wire \storeregister[14][5]~q ;
wire \storeregister[15][5]~feeder_combout ;
wire \storeregister[15][5]~q ;
wire \storeregister[13][5]~q ;
wire \storeregister[12][5]~q ;
wire \Mux26~17_combout ;
wire \Mux26~18_combout ;
wire \storeregister[5][5]~q ;
wire \storeregister[4][5]~q ;
wire \Mux26~10_combout ;
wire \storeregister[7][5]~q ;
wire \storeregister[6][5]~q ;
wire \Mux26~11_combout ;
wire \storeregister[24][3]~feeder_combout ;
wire \storeregister[24][3]~q ;
wire \Mux60~4_combout ;
wire \Mux60~5_combout ;
wire \Mux60~2_combout ;
wire \Mux60~3_combout ;
wire \Mux60~6_combout ;
wire \Mux60~0_combout ;
wire \Mux60~1_combout ;
wire \storeregister[19][3]~q ;
wire \Mux60~7_combout ;
wire \Mux60~8_combout ;
wire \Mux60~12_combout ;
wire \Mux60~13_combout ;
wire \storeregister[1][3]~q ;
wire \storeregister[3][3]~q ;
wire \Mux60~14_combout ;
wire \Mux60~15_combout ;
wire \Mux60~16_combout ;
wire \Mux60~17_combout ;
wire \Mux60~18_combout ;
wire \Mux60~10_combout ;
wire \Mux60~11_combout ;
wire \storeregister[29][16]~feeder_combout ;
wire \storeregister[29][16]~q ;
wire \storeregister[25][16]~feeder_combout ;
wire \storeregister[25][16]~q ;
wire \storeregister[17][16]~q ;
wire \storeregister[21][16]~q ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \storeregister[26][16]~feeder_combout ;
wire \storeregister[26][16]~q ;
wire \storeregister[18][16]~q ;
wire \Mux15~2_combout ;
wire \storeregister[30][16]~q ;
wire \storeregister[22][16]~feeder_combout ;
wire \storeregister[22][16]~q ;
wire \Mux15~3_combout ;
wire \storeregister[20][16]~q ;
wire \storeregister[16][16]~q ;
wire \storeregister[24][16]~feeder_combout ;
wire \storeregister[24][16]~q ;
wire \Mux15~4_combout ;
wire \Mux15~5_combout ;
wire \Mux15~6_combout ;
wire \storeregister[27][16]~feeder_combout ;
wire \storeregister[27][16]~q ;
wire \storeregister[23][16]~q ;
wire \Mux15~7_combout ;
wire \storeregister[31][16]~q ;
wire \Mux15~8_combout ;
wire \storeregister[10][16]~q ;
wire \storeregister[8][16]~feeder_combout ;
wire \storeregister[8][16]~q ;
wire \Mux15~10_combout ;
wire \storeregister[9][16]~q ;
wire \storeregister[11][16]~q ;
wire \Mux15~11_combout ;
wire \storeregister[4][16]~q ;
wire \storeregister[5][16]~q ;
wire \Mux15~12_combout ;
wire \storeregister[7][16]~q ;
wire \Mux15~13_combout ;
wire \storeregister[3][16]~q ;
wire \storeregister[1][16]~q ;
wire \Mux15~14_combout ;
wire \Mux15~15_combout ;
wire \Mux15~16_combout ;
wire \storeregister[14][16]~feeder_combout ;
wire \storeregister[14][16]~q ;
wire \storeregister[12][16]~q ;
wire \storeregister[13][16]~q ;
wire \Mux15~17_combout ;
wire \storeregister[15][16]~feeder_combout ;
wire \storeregister[15][16]~q ;
wire \Mux15~18_combout ;
wire \storeregister[31][14]~feeder_combout ;
wire \storeregister[31][14]~q ;
wire \storeregister[27][14]~q ;
wire \storeregister[19][14]~q ;
wire \storeregister[23][14]~q ;
wire \Mux17~7_combout ;
wire \Mux17~8_combout ;
wire \storeregister[30][14]~q ;
wire \storeregister[26][14]~feeder_combout ;
wire \storeregister[26][14]~q ;
wire \storeregister[18][14]~q ;
wire \Mux17~2_combout ;
wire \storeregister[22][14]~q ;
wire \Mux17~3_combout ;
wire \storeregister[16][14]~q ;
wire \storeregister[24][14]~q ;
wire \Mux17~4_combout ;
wire \storeregister[20][14]~q ;
wire \storeregister[28][14]~q ;
wire \Mux17~5_combout ;
wire \Mux17~6_combout ;
wire \storeregister[29][14]~feeder_combout ;
wire \storeregister[29][14]~q ;
wire \storeregister[25][14]~feeder_combout ;
wire \storeregister[25][14]~q ;
wire \storeregister[21][14]~feeder_combout ;
wire \storeregister[21][14]~q ;
wire \storeregister[17][14]~q ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \storeregister[12][14]~q ;
wire \storeregister[13][14]~feeder_combout ;
wire \storeregister[13][14]~q ;
wire \Mux17~17_combout ;
wire \storeregister[15][14]~feeder_combout ;
wire \storeregister[15][14]~q ;
wire \storeregister[14][14]~feeder_combout ;
wire \storeregister[14][14]~q ;
wire \Mux17~18_combout ;
wire \storeregister[9][14]~q ;
wire \storeregister[10][14]~q ;
wire \storeregister[8][14]~feeder_combout ;
wire \storeregister[8][14]~q ;
wire \Mux17~10_combout ;
wire \storeregister[11][14]~q ;
wire \Mux17~11_combout ;
wire \storeregister[6][14]~q ;
wire \storeregister[7][14]~q ;
wire \Mux17~13_combout ;
wire \storeregister[2][14]~q ;
wire \Mux17~15_combout ;
wire \Mux17~16_combout ;
wire \storeregister[28][15]~q ;
wire \storeregister[24][15]~q ;
wire \Mux16~5_combout ;
wire \storeregister[22][15]~q ;
wire \storeregister[18][15]~q ;
wire \Mux16~2_combout ;
wire \storeregister[30][15]~q ;
wire \storeregister[26][15]~feeder_combout ;
wire \storeregister[26][15]~q ;
wire \Mux16~3_combout ;
wire \Mux16~6_combout ;
wire \storeregister[29][15]~feeder_combout ;
wire \storeregister[29][15]~q ;
wire \storeregister[21][15]~q ;
wire \storeregister[25][15]~feeder_combout ;
wire \storeregister[25][15]~q ;
wire \storeregister[17][15]~q ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \storeregister[27][15]~q ;
wire \Mux16~7_combout ;
wire \storeregister[23][15]~feeder_combout ;
wire \storeregister[23][15]~q ;
wire \storeregister[31][15]~feeder_combout ;
wire \storeregister[31][15]~q ;
wire \Mux16~8_combout ;
wire \storeregister[7][15]~q ;
wire \storeregister[6][15]~q ;
wire \storeregister[4][15]~q ;
wire \storeregister[5][15]~q ;
wire \Mux16~10_combout ;
wire \Mux16~11_combout ;
wire \storeregister[15][15]~feeder_combout ;
wire \storeregister[15][15]~q ;
wire \storeregister[12][15]~q ;
wire \storeregister[13][15]~q ;
wire \Mux16~17_combout ;
wire \storeregister[14][15]~feeder_combout ;
wire \storeregister[14][15]~q ;
wire \Mux16~18_combout ;
wire \storeregister[3][15]~q ;
wire \storeregister[1][15]~q ;
wire \Mux16~14_combout ;
wire \storeregister[2][15]~q ;
wire \Mux16~15_combout ;
wire \storeregister[11][15]~q ;
wire \storeregister[9][15]~q ;
wire \Mux16~13_combout ;
wire \Mux16~16_combout ;
wire \storeregister[23][13]~q ;
wire \storeregister[27][13]~q ;
wire \storeregister[19][13]~q ;
wire \Mux18~7_combout ;
wire \storeregister[31][13]~q ;
wire \Mux18~8_combout ;
wire \storeregister[25][13]~q ;
wire \Mux18~0_combout ;
wire \storeregister[21][13]~feeder_combout ;
wire \storeregister[21][13]~q ;
wire \storeregister[29][13]~feeder_combout ;
wire \storeregister[29][13]~q ;
wire \Mux18~1_combout ;
wire \storeregister[22][13]~q ;
wire \storeregister[18][13]~q ;
wire \Mux18~2_combout ;
wire \storeregister[30][13]~q ;
wire \storeregister[26][13]~q ;
wire \Mux18~3_combout ;
wire \storeregister[24][13]~q ;
wire \storeregister[28][13]~feeder_combout ;
wire \storeregister[28][13]~q ;
wire \Mux18~5_combout ;
wire \Mux18~6_combout ;
wire \storeregister[11][13]~q ;
wire \storeregister[9][13]~q ;
wire \Mux18~13_combout ;
wire \storeregister[2][13]~feeder_combout ;
wire \storeregister[2][13]~q ;
wire \storeregister[1][13]~q ;
wire \storeregister[3][13]~q ;
wire \Mux18~14_combout ;
wire \Mux18~15_combout ;
wire \Mux18~16_combout ;
wire \storeregister[7][13]~q ;
wire \storeregister[6][13]~q ;
wire \storeregister[5][13]~q ;
wire \Mux18~10_combout ;
wire \Mux18~11_combout ;
wire \storeregister[14][13]~feeder_combout ;
wire \storeregister[14][13]~q ;
wire \storeregister[13][13]~q ;
wire \storeregister[12][13]~q ;
wire \Mux18~17_combout ;
wire \storeregister[15][13]~feeder_combout ;
wire \storeregister[15][13]~q ;
wire \Mux18~18_combout ;
wire \storeregister[29][12]~feeder_combout ;
wire \storeregister[29][12]~q ;
wire \storeregister[25][12]~q ;
wire \storeregister[17][12]~q ;
wire \storeregister[21][12]~q ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \storeregister[26][12]~q ;
wire \storeregister[18][12]~q ;
wire \Mux19~2_combout ;
wire \storeregister[22][12]~q ;
wire \storeregister[30][12]~feeder_combout ;
wire \storeregister[30][12]~q ;
wire \Mux19~3_combout ;
wire \storeregister[16][12]~q ;
wire \storeregister[24][12]~feeder_combout ;
wire \storeregister[24][12]~q ;
wire \Mux19~4_combout ;
wire \storeregister[28][12]~feeder_combout ;
wire \storeregister[28][12]~q ;
wire \storeregister[20][12]~q ;
wire \Mux19~5_combout ;
wire \Mux19~6_combout ;
wire \storeregister[19][12]~feeder_combout ;
wire \storeregister[19][12]~q ;
wire \storeregister[23][12]~q ;
wire \Mux19~7_combout ;
wire \storeregister[31][12]~feeder_combout ;
wire \storeregister[31][12]~q ;
wire \storeregister[27][12]~feeder_combout ;
wire \storeregister[27][12]~q ;
wire \Mux19~8_combout ;
wire \storeregister[7][12]~q ;
wire \storeregister[6][12]~q ;
wire \Mux19~13_combout ;
wire \storeregister[1][12]~q ;
wire \storeregister[3][12]~q ;
wire \Mux19~14_combout ;
wire \storeregister[2][12]~feeder_combout ;
wire \storeregister[2][12]~q ;
wire \Mux19~15_combout ;
wire \Mux19~16_combout ;
wire \storeregister[15][12]~feeder_combout ;
wire \storeregister[15][12]~q ;
wire \storeregister[14][12]~feeder_combout ;
wire \storeregister[14][12]~q ;
wire \storeregister[13][12]~q ;
wire \storeregister[12][12]~q ;
wire \Mux19~17_combout ;
wire \Mux19~18_combout ;
wire \storeregister[10][12]~q ;
wire \storeregister[8][12]~q ;
wire \Mux19~10_combout ;
wire \storeregister[9][12]~q ;
wire \storeregister[11][12]~q ;
wire \Mux19~11_combout ;
wire \storeregister[28][10]~q ;
wire \storeregister[20][10]~q ;
wire \Mux21~5_combout ;
wire \storeregister[26][10]~q ;
wire \Mux21~2_combout ;
wire \storeregister[22][10]~q ;
wire \storeregister[30][10]~q ;
wire \Mux21~3_combout ;
wire \Mux21~6_combout ;
wire \storeregister[21][10]~feeder_combout ;
wire \storeregister[21][10]~q ;
wire \storeregister[17][10]~q ;
wire \Mux21~0_combout ;
wire \storeregister[25][10]~q ;
wire \storeregister[29][10]~q ;
wire \Mux21~1_combout ;
wire \storeregister[19][10]~q ;
wire \storeregister[23][10]~q ;
wire \Mux21~7_combout ;
wire \storeregister[27][10]~q ;
wire \storeregister[31][10]~feeder_combout ;
wire \storeregister[31][10]~q ;
wire \Mux21~8_combout ;
wire \storeregister[8][10]~feeder_combout ;
wire \storeregister[8][10]~q ;
wire \storeregister[10][10]~q ;
wire \Mux21~10_combout ;
wire \storeregister[9][10]~q ;
wire \storeregister[11][10]~q ;
wire \Mux21~11_combout ;
wire \storeregister[7][10]~q ;
wire \storeregister[4][10]~q ;
wire \storeregister[5][10]~q ;
wire \Mux21~12_combout ;
wire \Mux21~13_combout ;
wire \storeregister[2][10]~feeder_combout ;
wire \storeregister[2][10]~q ;
wire \storeregister[3][10]~q ;
wire \Mux21~14_combout ;
wire \Mux21~15_combout ;
wire \Mux21~16_combout ;
wire \storeregister[12][10]~q ;
wire \storeregister[13][10]~q ;
wire \Mux21~17_combout ;
wire \storeregister[14][10]~feeder_combout ;
wire \storeregister[14][10]~q ;
wire \storeregister[15][10]~q ;
wire \Mux21~18_combout ;
wire \storeregister[26][11]~q ;
wire \storeregister[22][11]~q ;
wire \storeregister[18][11]~q ;
wire \Mux20~2_combout ;
wire \Mux20~3_combout ;
wire \storeregister[28][11]~feeder_combout ;
wire \storeregister[28][11]~q ;
wire \storeregister[16][11]~q ;
wire \Mux20~4_combout ;
wire \Mux20~5_combout ;
wire \Mux20~6_combout ;
wire \storeregister[21][11]~feeder_combout ;
wire \storeregister[21][11]~q ;
wire \storeregister[29][11]~feeder_combout ;
wire \storeregister[29][11]~q ;
wire \storeregister[25][11]~q ;
wire \storeregister[17][11]~feeder_combout ;
wire \storeregister[17][11]~q ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \storeregister[31][11]~feeder_combout ;
wire \storeregister[31][11]~q ;
wire \storeregister[19][11]~feeder_combout ;
wire \storeregister[19][11]~q ;
wire \Mux20~7_combout ;
wire \storeregister[23][11]~q ;
wire \Mux20~8_combout ;
wire \storeregister[7][11]~feeder_combout ;
wire \storeregister[7][11]~q ;
wire \storeregister[5][11]~q ;
wire \storeregister[4][11]~q ;
wire \Mux20~10_combout ;
wire \storeregister[6][11]~feeder_combout ;
wire \storeregister[6][11]~q ;
wire \Mux20~11_combout ;
wire \storeregister[3][11]~q ;
wire \Mux20~14_combout ;
wire \storeregister[2][11]~q ;
wire \Mux20~15_combout ;
wire \storeregister[11][11]~feeder_combout ;
wire \storeregister[11][11]~q ;
wire \storeregister[9][11]~feeder_combout ;
wire \storeregister[9][11]~q ;
wire \Mux20~13_combout ;
wire \Mux20~16_combout ;
wire \storeregister[15][11]~feeder_combout ;
wire \storeregister[15][11]~q ;
wire \storeregister[14][11]~feeder_combout ;
wire \storeregister[14][11]~q ;
wire \storeregister[13][11]~q ;
wire \storeregister[12][11]~q ;
wire \Mux20~17_combout ;
wire \Mux20~18_combout ;
wire \storeregister[17][9]~q ;
wire \Mux22~0_combout ;
wire \storeregister[29][9]~feeder_combout ;
wire \storeregister[29][9]~q ;
wire \storeregister[21][9]~feeder_combout ;
wire \storeregister[21][9]~q ;
wire \Mux22~1_combout ;
wire \storeregister[30][9]~q ;
wire \storeregister[26][9]~q ;
wire \Mux22~3_combout ;
wire \storeregister[28][9]~q ;
wire \storeregister[24][9]~feeder_combout ;
wire \storeregister[24][9]~q ;
wire \Mux22~5_combout ;
wire \Mux22~6_combout ;
wire \storeregister[23][9]~q ;
wire \storeregister[31][9]~q ;
wire \storeregister[19][9]~q ;
wire \storeregister[27][9]~feeder_combout ;
wire \storeregister[27][9]~q ;
wire \Mux22~7_combout ;
wire \Mux22~8_combout ;
wire \storeregister[5][9]~q ;
wire \Mux22~10_combout ;
wire \storeregister[7][9]~q ;
wire \storeregister[6][9]~q ;
wire \Mux22~11_combout ;
wire \storeregister[12][9]~q ;
wire \storeregister[13][9]~q ;
wire \Mux22~17_combout ;
wire \storeregister[14][9]~q ;
wire \storeregister[15][9]~feeder_combout ;
wire \storeregister[15][9]~q ;
wire \Mux22~18_combout ;
wire \storeregister[8][9]~q ;
wire \storeregister[10][9]~q ;
wire \Mux22~12_combout ;
wire \storeregister[11][9]~q ;
wire \storeregister[9][9]~q ;
wire \Mux22~13_combout ;
wire \storeregister[2][9]~q ;
wire \storeregister[3][9]~q ;
wire \Mux22~14_combout ;
wire \Mux22~15_combout ;
wire \Mux22~16_combout ;
wire \Mux59~7_combout ;
wire \Mux59~8_combout ;
wire \Mux59~0_combout ;
wire \Mux59~1_combout ;
wire \Mux59~5_combout ;
wire \Mux59~3_combout ;
wire \Mux59~6_combout ;
wire \Mux59~13_combout ;
wire \Mux59~14_combout ;
wire \storeregister[2][4]~q ;
wire \Mux59~15_combout ;
wire \Mux59~16_combout ;
wire \Mux59~17_combout ;
wire \Mux59~18_combout ;
wire \Mux59~10_combout ;
wire \storeregister[6][4]~feeder_combout ;
wire \storeregister[6][4]~q ;
wire \Mux59~11_combout ;
wire \storeregister[27][31]~feeder_combout ;
wire \storeregister[27][31]~q ;
wire \storeregister[19][31]~q ;
wire \Mux0~7_combout ;
wire \storeregister[31][31]~q ;
wire \storeregister[23][31]~feeder_combout ;
wire \storeregister[23][31]~q ;
wire \Mux0~8_combout ;
wire \storeregister[26][31]~feeder_combout ;
wire \storeregister[26][31]~q ;
wire \storeregister[30][31]~feeder_combout ;
wire \storeregister[30][31]~q ;
wire \Mux0~3_combout ;
wire \storeregister[20][31]~q ;
wire \Mux0~4_combout ;
wire \storeregister[24][31]~feeder_combout ;
wire \storeregister[24][31]~q ;
wire \Mux0~5_combout ;
wire \Mux0~6_combout ;
wire \storeregister[25][31]~q ;
wire \Mux0~0_combout ;
wire \storeregister[21][31]~q ;
wire \storeregister[29][31]~q ;
wire \Mux0~1_combout ;
wire \storeregister[15][31]~feeder_combout ;
wire \storeregister[15][31]~q ;
wire \storeregister[14][31]~q ;
wire \storeregister[12][31]~q ;
wire \Mux0~17_combout ;
wire \Mux0~18_combout ;
wire \storeregister[2][31]~q ;
wire \storeregister[3][31]~q ;
wire \Mux0~14_combout ;
wire \Mux0~15_combout ;
wire \storeregister[9][31]~feeder_combout ;
wire \storeregister[9][31]~q ;
wire \storeregister[11][31]~q ;
wire \Mux0~13_combout ;
wire \Mux0~16_combout ;
wire \storeregister[5][31]~q ;
wire \storeregister[4][31]~q ;
wire \Mux0~10_combout ;
wire \storeregister[6][31]~q ;
wire \storeregister[7][31]~q ;
wire \Mux0~11_combout ;
wire \storeregister[29][30]~q ;
wire \storeregister[21][30]~q ;
wire \storeregister[17][30]~feeder_combout ;
wire \storeregister[17][30]~q ;
wire \Mux1~0_combout ;
wire \storeregister[25][30]~q ;
wire \Mux1~1_combout ;
wire \storeregister[30][30]~q ;
wire \storeregister[26][30]~q ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \storeregister[20][30]~q ;
wire \storeregister[28][30]~q ;
wire \storeregister[16][30]~q ;
wire \storeregister[24][30]~q ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux1~6_combout ;
wire \storeregister[23][30]~q ;
wire \storeregister[19][30]~q ;
wire \Mux1~7_combout ;
wire \storeregister[31][30]~q ;
wire \storeregister[27][30]~q ;
wire \Mux1~8_combout ;
wire \storeregister[15][30]~feeder_combout ;
wire \storeregister[15][30]~q ;
wire \storeregister[14][30]~feeder_combout ;
wire \storeregister[14][30]~q ;
wire \storeregister[13][30]~q ;
wire \storeregister[12][30]~q ;
wire \Mux1~17_combout ;
wire \Mux1~18_combout ;
wire \storeregister[7][30]~q ;
wire \storeregister[6][30]~q ;
wire \Mux1~13_combout ;
wire \storeregister[2][30]~q ;
wire \storeregister[1][30]~q ;
wire \storeregister[3][30]~q ;
wire \Mux1~14_combout ;
wire \Mux1~15_combout ;
wire \Mux1~16_combout ;
wire \storeregister[10][30]~q ;
wire \Mux1~10_combout ;
wire \storeregister[11][30]~q ;
wire \storeregister[9][30]~q ;
wire \Mux1~11_combout ;
wire \storeregister[30][29]~q ;
wire \storeregister[26][29]~q ;
wire \storeregister[22][29]~q ;
wire \storeregister[18][29]~q ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;
wire \storeregister[24][29]~q ;
wire \storeregister[16][29]~q ;
wire \Mux2~4_combout ;
wire \Mux2~5_combout ;
wire \Mux2~6_combout ;
wire \storeregister[29][29]~feeder_combout ;
wire \storeregister[29][29]~q ;
wire \storeregister[25][29]~q ;
wire \storeregister[17][29]~q ;
wire \Mux2~0_combout ;
wire \storeregister[21][29]~feeder_combout ;
wire \storeregister[21][29]~q ;
wire \Mux2~1_combout ;
wire \storeregister[27][29]~q ;
wire \storeregister[19][29]~q ;
wire \Mux2~7_combout ;
wire \storeregister[31][29]~q ;
wire \storeregister[23][29]~feeder_combout ;
wire \storeregister[23][29]~q ;
wire \Mux2~8_combout ;
wire \storeregister[12][29]~feeder_combout ;
wire \storeregister[12][29]~q ;
wire \storeregister[13][29]~q ;
wire \Mux2~17_combout ;
wire \storeregister[14][29]~q ;
wire \storeregister[15][29]~feeder_combout ;
wire \storeregister[15][29]~q ;
wire \Mux2~18_combout ;
wire \storeregister[9][29]~feeder_combout ;
wire \storeregister[9][29]~q ;
wire \storeregister[11][29]~q ;
wire \storeregister[10][29]~q ;
wire \storeregister[8][29]~q ;
wire \Mux2~12_combout ;
wire \Mux2~13_combout ;
wire \storeregister[2][29]~q ;
wire \Mux2~15_combout ;
wire \Mux2~16_combout ;
wire \storeregister[7][29]~q ;
wire \storeregister[6][29]~q ;
wire \storeregister[5][29]~q ;
wire \storeregister[4][29]~q ;
wire \Mux2~10_combout ;
wire \Mux2~11_combout ;
wire \storeregister[23][26]~feeder_combout ;
wire \storeregister[23][26]~q ;
wire \storeregister[19][26]~q ;
wire \Mux5~7_combout ;
wire \storeregister[31][26]~q ;
wire \storeregister[27][26]~q ;
wire \Mux5~8_combout ;
wire \storeregister[16][26]~q ;
wire \storeregister[24][26]~q ;
wire \Mux5~4_combout ;
wire \storeregister[28][26]~feeder_combout ;
wire \storeregister[28][26]~q ;
wire \Mux5~5_combout ;
wire \storeregister[26][26]~q ;
wire \Mux5~2_combout ;
wire \storeregister[22][26]~q ;
wire \storeregister[30][26]~feeder_combout ;
wire \storeregister[30][26]~q ;
wire \Mux5~3_combout ;
wire \Mux5~6_combout ;
wire \storeregister[29][26]~feeder_combout ;
wire \storeregister[29][26]~q ;
wire \storeregister[21][26]~feeder_combout ;
wire \storeregister[21][26]~q ;
wire \Mux5~0_combout ;
wire \storeregister[25][26]~q ;
wire \Mux5~1_combout ;
wire \storeregister[9][26]~feeder_combout ;
wire \storeregister[9][26]~q ;
wire \storeregister[11][26]~q ;
wire \storeregister[10][26]~q ;
wire \Mux5~10_combout ;
wire \Mux5~11_combout ;
wire \storeregister[14][26]~q ;
wire \storeregister[15][26]~feeder_combout ;
wire \storeregister[15][26]~q ;
wire \storeregister[13][26]~q ;
wire \storeregister[12][26]~q ;
wire \Mux5~17_combout ;
wire \Mux5~18_combout ;
wire \storeregister[2][26]~q ;
wire \storeregister[3][26]~q ;
wire \Mux5~14_combout ;
wire \Mux5~15_combout ;
wire \storeregister[7][26]~q ;
wire \storeregister[6][26]~q ;
wire \Mux5~13_combout ;
wire \Mux5~16_combout ;
wire \storeregister[30][25]~feeder_combout ;
wire \storeregister[30][25]~q ;
wire \storeregister[18][25]~q ;
wire \storeregister[22][25]~q ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \storeregister[16][25]~q ;
wire \storeregister[20][25]~feeder_combout ;
wire \storeregister[20][25]~q ;
wire \Mux6~4_combout ;
wire \storeregister[28][25]~q ;
wire \Mux6~5_combout ;
wire \Mux6~6_combout ;
wire \storeregister[31][25]~q ;
wire \storeregister[19][25]~feeder_combout ;
wire \storeregister[19][25]~q ;
wire \storeregister[27][25]~q ;
wire \Mux6~7_combout ;
wire \storeregister[23][25]~q ;
wire \Mux6~8_combout ;
wire \storeregister[29][25]~feeder_combout ;
wire \storeregister[29][25]~q ;
wire \storeregister[21][25]~feeder_combout ;
wire \storeregister[21][25]~q ;
wire \storeregister[25][25]~q ;
wire \storeregister[17][25]~feeder_combout ;
wire \storeregister[17][25]~q ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \storeregister[15][25]~feeder_combout ;
wire \storeregister[15][25]~q ;
wire \storeregister[12][25]~q ;
wire \storeregister[13][25]~q ;
wire \Mux6~17_combout ;
wire \storeregister[14][25]~q ;
wire \Mux6~18_combout ;
wire \storeregister[9][25]~q ;
wire \storeregister[11][25]~q ;
wire \Mux6~13_combout ;
wire \storeregister[2][25]~q ;
wire \storeregister[3][25]~q ;
wire \Mux6~14_combout ;
wire \Mux6~15_combout ;
wire \Mux6~16_combout ;
wire \storeregister[7][25]~q ;
wire \storeregister[6][25]~q ;
wire \storeregister[5][25]~q ;
wire \Mux6~10_combout ;
wire \Mux6~11_combout ;
wire \storeregister[20][28]~q ;
wire \storeregister[16][28]~feeder_combout ;
wire \storeregister[16][28]~q ;
wire \storeregister[24][28]~feeder_combout ;
wire \storeregister[24][28]~q ;
wire \Mux3~4_combout ;
wire \Mux3~5_combout ;
wire \storeregister[30][28]~feeder_combout ;
wire \storeregister[30][28]~q ;
wire \storeregister[26][28]~q ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \Mux3~6_combout ;
wire \storeregister[31][28]~q ;
wire \storeregister[19][28]~feeder_combout ;
wire \storeregister[19][28]~q ;
wire \storeregister[23][28]~q ;
wire \Mux3~7_combout ;
wire \storeregister[27][28]~q ;
wire \Mux3~8_combout ;
wire \storeregister[25][28]~q ;
wire \storeregister[29][28]~q ;
wire \storeregister[21][28]~feeder_combout ;
wire \storeregister[21][28]~q ;
wire \storeregister[17][28]~q ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \storeregister[10][28]~q ;
wire \Mux3~10_combout ;
wire \storeregister[9][28]~q ;
wire \storeregister[11][28]~q ;
wire \Mux3~11_combout ;
wire \storeregister[15][28]~q ;
wire \storeregister[12][28]~feeder_combout ;
wire \storeregister[12][28]~q ;
wire \storeregister[13][28]~feeder_combout ;
wire \storeregister[13][28]~q ;
wire \Mux3~17_combout ;
wire \storeregister[14][28]~feeder_combout ;
wire \storeregister[14][28]~q ;
wire \Mux3~18_combout ;
wire \storeregister[2][28]~q ;
wire \storeregister[3][28]~q ;
wire \Mux3~14_combout ;
wire \Mux3~15_combout ;
wire \storeregister[7][28]~q ;
wire \storeregister[6][28]~q ;
wire \Mux3~13_combout ;
wire \Mux3~16_combout ;
wire \storeregister[27][27]~q ;
wire \storeregister[19][27]~q ;
wire \Mux4~7_combout ;
wire \storeregister[23][27]~q ;
wire \storeregister[31][27]~feeder_combout ;
wire \storeregister[31][27]~q ;
wire \Mux4~8_combout ;
wire \storeregister[25][27]~q ;
wire \storeregister[17][27]~q ;
wire \Mux4~0_combout ;
wire \storeregister[29][27]~q ;
wire \storeregister[21][27]~feeder_combout ;
wire \storeregister[21][27]~q ;
wire \Mux4~1_combout ;
wire \storeregister[26][27]~q ;
wire \storeregister[30][27]~q ;
wire \Mux4~3_combout ;
wire \storeregister[20][27]~q ;
wire \storeregister[16][27]~q ;
wire \Mux4~4_combout ;
wire \storeregister[28][27]~q ;
wire \Mux4~5_combout ;
wire \Mux4~6_combout ;
wire \storeregister[6][27]~q ;
wire \storeregister[7][27]~q ;
wire \storeregister[5][27]~q ;
wire \storeregister[4][27]~q ;
wire \Mux4~10_combout ;
wire \Mux4~11_combout ;
wire \storeregister[10][27]~q ;
wire \storeregister[8][27]~q ;
wire \Mux4~12_combout ;
wire \storeregister[11][27]~q ;
wire \Mux4~13_combout ;
wire \storeregister[1][27]~q ;
wire \storeregister[3][27]~q ;
wire \Mux4~14_combout ;
wire \storeregister[2][27]~q ;
wire \Mux4~15_combout ;
wire \Mux4~16_combout ;
wire \storeregister[15][27]~feeder_combout ;
wire \storeregister[15][27]~q ;
wire \storeregister[14][27]~feeder_combout ;
wire \storeregister[14][27]~q ;
wire \storeregister[12][27]~q ;
wire \Mux4~17_combout ;
wire \Mux4~18_combout ;
wire \storeregister[26][17]~feeder_combout ;
wire \storeregister[26][17]~q ;
wire \storeregister[30][17]~feeder_combout ;
wire \storeregister[30][17]~q ;
wire \Mux14~3_combout ;
wire \storeregister[16][17]~q ;
wire \Mux14~4_combout ;
wire \storeregister[24][17]~q ;
wire \Mux14~5_combout ;
wire \Mux14~6_combout ;
wire \storeregister[23][17]~q ;
wire \storeregister[31][17]~q ;
wire \storeregister[27][17]~feeder_combout ;
wire \storeregister[27][17]~q ;
wire \storeregister[19][17]~q ;
wire \Mux14~7_combout ;
wire \Mux14~8_combout ;
wire \storeregister[21][17]~q ;
wire \storeregister[25][17]~q ;
wire \storeregister[17][17]~q ;
wire \Mux14~0_combout ;
wire \storeregister[29][17]~q ;
wire \Mux14~1_combout ;
wire \storeregister[14][17]~feeder_combout ;
wire \storeregister[14][17]~q ;
wire \storeregister[12][17]~q ;
wire \storeregister[13][17]~q ;
wire \Mux14~17_combout ;
wire \storeregister[15][17]~feeder_combout ;
wire \storeregister[15][17]~q ;
wire \Mux14~18_combout ;
wire \storeregister[2][17]~q ;
wire \storeregister[1][17]~q ;
wire \storeregister[3][17]~q ;
wire \Mux14~14_combout ;
wire \Mux14~15_combout ;
wire \storeregister[8][17]~q ;
wire \storeregister[10][17]~q ;
wire \Mux14~12_combout ;
wire \storeregister[11][17]~q ;
wire \Mux14~13_combout ;
wire \Mux14~16_combout ;
wire \storeregister[5][17]~q ;
wire \storeregister[4][17]~q ;
wire \Mux14~10_combout ;
wire \storeregister[6][17]~q ;
wire \storeregister[7][17]~q ;
wire \Mux14~11_combout ;
wire \storeregister[31][20]~q ;
wire \storeregister[27][20]~q ;
wire \storeregister[19][20]~q ;
wire \Mux11~7_combout ;
wire \Mux11~8_combout ;
wire \storeregister[25][20]~q ;
wire \storeregister[29][20]~q ;
wire \storeregister[21][20]~feeder_combout ;
wire \storeregister[21][20]~q ;
wire \storeregister[17][20]~q ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \storeregister[20][20]~q ;
wire \storeregister[28][20]~q ;
wire \Mux11~5_combout ;
wire \storeregister[30][20]~q ;
wire \storeregister[22][20]~q ;
wire \storeregister[26][20]~feeder_combout ;
wire \storeregister[26][20]~q ;
wire \storeregister[18][20]~q ;
wire \Mux11~2_combout ;
wire \Mux11~3_combout ;
wire \Mux11~6_combout ;
wire \storeregister[15][20]~feeder_combout ;
wire \storeregister[15][20]~q ;
wire \storeregister[12][20]~q ;
wire \storeregister[13][20]~q ;
wire \Mux11~17_combout ;
wire \storeregister[14][20]~feeder_combout ;
wire \storeregister[14][20]~q ;
wire \Mux11~18_combout ;
wire \storeregister[2][20]~q ;
wire \Mux11~15_combout ;
wire \storeregister[6][20]~q ;
wire \storeregister[7][20]~q ;
wire \storeregister[5][20]~q ;
wire \storeregister[4][20]~q ;
wire \Mux11~12_combout ;
wire \Mux11~13_combout ;
wire \Mux11~16_combout ;
wire \storeregister[8][20]~q ;
wire \storeregister[10][20]~q ;
wire \Mux11~10_combout ;
wire \storeregister[9][20]~q ;
wire \storeregister[11][20]~q ;
wire \Mux11~11_combout ;
wire \storeregister[30][19]~q ;
wire \storeregister[22][19]~q ;
wire \storeregister[18][19]~q ;
wire \Mux12~2_combout ;
wire \Mux12~3_combout ;
wire \storeregister[28][19]~q ;
wire \storeregister[16][19]~q ;
wire \storeregister[20][19]~q ;
wire \Mux12~4_combout ;
wire \Mux12~5_combout ;
wire \Mux12~6_combout ;
wire \storeregister[25][19]~q ;
wire \storeregister[17][19]~q ;
wire \Mux12~0_combout ;
wire \storeregister[29][19]~q ;
wire \storeregister[21][19]~q ;
wire \Mux12~1_combout ;
wire \storeregister[19][19]~feeder_combout ;
wire \storeregister[19][19]~q ;
wire \storeregister[27][19]~feeder_combout ;
wire \storeregister[27][19]~q ;
wire \Mux12~7_combout ;
wire \storeregister[31][19]~feeder_combout ;
wire \storeregister[31][19]~q ;
wire \storeregister[23][19]~feeder_combout ;
wire \storeregister[23][19]~q ;
wire \Mux12~8_combout ;
wire \storeregister[14][19]~feeder_combout ;
wire \storeregister[14][19]~q ;
wire \storeregister[15][19]~feeder_combout ;
wire \storeregister[15][19]~q ;
wire \storeregister[13][19]~q ;
wire \storeregister[12][19]~q ;
wire \Mux12~17_combout ;
wire \Mux12~18_combout ;
wire \storeregister[9][19]~q ;
wire \storeregister[11][19]~q ;
wire \Mux12~13_combout ;
wire \storeregister[2][19]~q ;
wire \storeregister[1][19]~q ;
wire \storeregister[3][19]~q ;
wire \Mux12~14_combout ;
wire \Mux12~15_combout ;
wire \Mux12~16_combout ;
wire \storeregister[6][19]~feeder_combout ;
wire \storeregister[6][19]~q ;
wire \storeregister[5][19]~q ;
wire \Mux12~10_combout ;
wire \storeregister[7][19]~q ;
wire \Mux12~11_combout ;
wire \storeregister[28][18]~feeder_combout ;
wire \storeregister[28][18]~q ;
wire \storeregister[20][18]~feeder_combout ;
wire \storeregister[20][18]~q ;
wire \storeregister[24][18]~q ;
wire \Mux13~4_combout ;
wire \Mux13~5_combout ;
wire \storeregister[30][18]~q ;
wire \storeregister[22][18]~feeder_combout ;
wire \storeregister[22][18]~q ;
wire \Mux13~3_combout ;
wire \Mux13~6_combout ;
wire \storeregister[27][18]~q ;
wire \storeregister[31][18]~q ;
wire \storeregister[23][18]~q ;
wire \storeregister[19][18]~q ;
wire \Mux13~7_combout ;
wire \Mux13~8_combout ;
wire \storeregister[29][18]~q ;
wire \storeregister[17][18]~feeder_combout ;
wire \storeregister[17][18]~q ;
wire \storeregister[21][18]~q ;
wire \Mux13~0_combout ;
wire \storeregister[25][18]~q ;
wire \Mux13~1_combout ;
wire \storeregister[15][18]~feeder_combout ;
wire \storeregister[15][18]~q ;
wire \storeregister[14][18]~feeder_combout ;
wire \storeregister[14][18]~q ;
wire \storeregister[13][18]~q ;
wire \storeregister[12][18]~q ;
wire \Mux13~17_combout ;
wire \Mux13~18_combout ;
wire \storeregister[11][18]~q ;
wire \storeregister[10][18]~q ;
wire \storeregister[8][18]~q ;
wire \Mux13~10_combout ;
wire \storeregister[9][18]~q ;
wire \Mux13~11_combout ;
wire \storeregister[2][18]~feeder_combout ;
wire \storeregister[2][18]~q ;
wire \Mux13~15_combout ;
wire \storeregister[4][18]~q ;
wire \storeregister[5][18]~q ;
wire \Mux13~12_combout ;
wire \storeregister[7][18]~q ;
wire \storeregister[6][18]~q ;
wire \Mux13~13_combout ;
wire \Mux13~16_combout ;
wire \storeregister[29][24]~q ;
wire \storeregister[25][24]~q ;
wire \storeregister[21][24]~q ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \storeregister[19][24]~q ;
wire \Mux7~7_combout ;
wire \storeregister[31][24]~feeder_combout ;
wire \storeregister[31][24]~q ;
wire \storeregister[27][24]~q ;
wire \Mux7~8_combout ;
wire \storeregister[30][24]~feeder_combout ;
wire \storeregister[30][24]~q ;
wire \storeregister[26][24]~q ;
wire \storeregister[18][24]~q ;
wire \Mux7~2_combout ;
wire \Mux7~3_combout ;
wire \storeregister[28][24]~feeder_combout ;
wire \storeregister[28][24]~q ;
wire \storeregister[16][24]~q ;
wire \storeregister[24][24]~feeder_combout ;
wire \storeregister[24][24]~q ;
wire \Mux7~4_combout ;
wire \Mux7~5_combout ;
wire \Mux7~6_combout ;
wire \storeregister[13][24]~q ;
wire \Mux7~17_combout ;
wire \storeregister[14][24]~feeder_combout ;
wire \storeregister[14][24]~q ;
wire \storeregister[15][24]~feeder_combout ;
wire \storeregister[15][24]~q ;
wire \Mux7~18_combout ;
wire \storeregister[10][24]~q ;
wire \storeregister[8][24]~q ;
wire \Mux7~10_combout ;
wire \storeregister[9][24]~q ;
wire \storeregister[11][24]~q ;
wire \Mux7~11_combout ;
wire \storeregister[4][24]~q ;
wire \Mux7~12_combout ;
wire \storeregister[7][24]~q ;
wire \Mux7~13_combout ;
wire \storeregister[2][24]~feeder_combout ;
wire \storeregister[2][24]~q ;
wire \storeregister[3][24]~q ;
wire \Mux7~14_combout ;
wire \Mux7~15_combout ;
wire \Mux7~16_combout ;
wire \storeregister[30][23]~q ;
wire \storeregister[26][23]~q ;
wire \Mux8~3_combout ;
wire \storeregister[28][23]~feeder_combout ;
wire \storeregister[28][23]~q ;
wire \storeregister[24][23]~q ;
wire \storeregister[16][23]~q ;
wire \storeregister[20][23]~q ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \Mux8~6_combout ;
wire \storeregister[21][23]~feeder_combout ;
wire \storeregister[21][23]~q ;
wire \storeregister[29][23]~q ;
wire \storeregister[25][23]~q ;
wire \storeregister[17][23]~q ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \storeregister[23][23]~q ;
wire \storeregister[19][23]~feeder_combout ;
wire \storeregister[19][23]~q ;
wire \storeregister[27][23]~q ;
wire \Mux8~7_combout ;
wire \storeregister[31][23]~q ;
wire \Mux8~8_combout ;
wire \storeregister[5][23]~q ;
wire \storeregister[4][23]~q ;
wire \Mux8~10_combout ;
wire \storeregister[6][23]~q ;
wire \storeregister[7][23]~q ;
wire \Mux8~11_combout ;
wire \storeregister[2][23]~feeder_combout ;
wire \storeregister[2][23]~q ;
wire \storeregister[3][23]~q ;
wire \storeregister[1][23]~q ;
wire \Mux8~14_combout ;
wire \Mux8~15_combout ;
wire \storeregister[11][23]~q ;
wire \storeregister[9][23]~q ;
wire \Mux8~13_combout ;
wire \Mux8~16_combout ;
wire \storeregister[13][23]~q ;
wire \storeregister[12][23]~q ;
wire \Mux8~17_combout ;
wire \storeregister[14][23]~feeder_combout ;
wire \storeregister[14][23]~q ;
wire \storeregister[15][23]~feeder_combout ;
wire \storeregister[15][23]~q ;
wire \Mux8~18_combout ;
wire \storeregister[27][22]~q ;
wire \storeregister[19][22]~q ;
wire \storeregister[23][22]~feeder_combout ;
wire \storeregister[23][22]~q ;
wire \Mux9~7_combout ;
wire \storeregister[31][22]~q ;
wire \Mux9~8_combout ;
wire \storeregister[25][22]~q ;
wire \storeregister[17][22]~q ;
wire \Mux9~0_combout ;
wire \storeregister[29][22]~q ;
wire \Mux9~1_combout ;
wire \storeregister[30][22]~q ;
wire \storeregister[22][22]~q ;
wire \Mux9~3_combout ;
wire \storeregister[28][22]~q ;
wire \storeregister[16][22]~q ;
wire \storeregister[24][22]~feeder_combout ;
wire \storeregister[24][22]~q ;
wire \Mux9~4_combout ;
wire \Mux9~5_combout ;
wire \Mux9~6_combout ;
wire \storeregister[10][22]~q ;
wire \Mux9~10_combout ;
wire \storeregister[9][22]~q ;
wire \storeregister[11][22]~q ;
wire \Mux9~11_combout ;
wire \storeregister[14][22]~feeder_combout ;
wire \storeregister[14][22]~q ;
wire \storeregister[15][22]~q ;
wire \storeregister[13][22]~q ;
wire \storeregister[12][22]~q ;
wire \Mux9~17_combout ;
wire \Mux9~18_combout ;
wire \storeregister[4][22]~q ;
wire \storeregister[5][22]~q ;
wire \Mux9~12_combout ;
wire \storeregister[7][22]~q ;
wire \storeregister[6][22]~q ;
wire \Mux9~13_combout ;
wire \storeregister[2][22]~q ;
wire \Mux9~15_combout ;
wire \Mux9~16_combout ;
wire \storeregister[24][21]~feeder_combout ;
wire \storeregister[24][21]~q ;
wire \storeregister[28][21]~q ;
wire \Mux10~5_combout ;
wire \storeregister[22][21]~q ;
wire \storeregister[18][21]~q ;
wire \Mux10~2_combout ;
wire \storeregister[26][21]~q ;
wire \Mux10~3_combout ;
wire \Mux10~6_combout ;
wire \storeregister[21][21]~q ;
wire \storeregister[29][21]~q ;
wire \storeregister[25][21]~feeder_combout ;
wire \storeregister[25][21]~q ;
wire \storeregister[17][21]~q ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \storeregister[27][21]~feeder_combout ;
wire \storeregister[27][21]~q ;
wire \storeregister[19][21]~feeder_combout ;
wire \storeregister[19][21]~q ;
wire \Mux10~7_combout ;
wire \storeregister[31][21]~q ;
wire \storeregister[23][21]~q ;
wire \Mux10~8_combout ;
wire \storeregister[8][21]~q ;
wire \storeregister[10][21]~q ;
wire \Mux10~12_combout ;
wire \storeregister[11][21]~q ;
wire \Mux10~13_combout ;
wire \storeregister[3][21]~q ;
wire \storeregister[1][21]~q ;
wire \Mux10~14_combout ;
wire \Mux10~15_combout ;
wire \Mux10~16_combout ;
wire \storeregister[15][21]~feeder_combout ;
wire \storeregister[15][21]~q ;
wire \storeregister[13][21]~q ;
wire \storeregister[12][21]~q ;
wire \Mux10~17_combout ;
wire \storeregister[14][21]~feeder_combout ;
wire \storeregister[14][21]~q ;
wire \Mux10~18_combout ;
wire \storeregister[7][21]~q ;
wire \storeregister[6][21]~q ;
wire \storeregister[5][21]~q ;
wire \storeregister[4][21]~q ;
wire \Mux10~10_combout ;
wire \Mux10~11_combout ;
wire \storeregister[20][15]~q ;
wire \storeregister[16][15]~q ;
wire \Mux48~4_combout ;
wire \Mux48~5_combout ;
wire \Mux48~3_combout ;
wire \Mux48~6_combout ;
wire \storeregister[19][15]~feeder_combout ;
wire \storeregister[19][15]~q ;
wire \Mux48~7_combout ;
wire \Mux48~8_combout ;
wire \Mux48~0_combout ;
wire \Mux48~1_combout ;
wire \Mux48~17_combout ;
wire \Mux48~18_combout ;
wire \Mux48~12_combout ;
wire \Mux48~13_combout ;
wire \Mux48~14_combout ;
wire \Mux48~15_combout ;
wire \Mux48~16_combout ;
wire \storeregister[10][15]~q ;
wire \storeregister[8][15]~q ;
wire \Mux48~10_combout ;
wire \Mux48~11_combout ;
wire \Mux51~7_combout ;
wire \Mux51~8_combout ;
wire \Mux51~0_combout ;
wire \Mux51~1_combout ;
wire \Mux51~2_combout ;
wire \Mux51~3_combout ;
wire \Mux51~4_combout ;
wire \Mux51~5_combout ;
wire \Mux51~6_combout ;
wire \Mux51~12_combout ;
wire \Mux51~13_combout ;
wire \Mux51~14_combout ;
wire \Mux51~15_combout ;
wire \Mux51~16_combout ;
wire \Mux51~17_combout ;
wire \Mux51~18_combout ;
wire \storeregister[4][12]~q ;
wire \storeregister[5][12]~q ;
wire \Mux51~10_combout ;
wire \Mux51~11_combout ;
wire \storeregister[22][27]~q ;
wire \storeregister[18][27]~q ;
wire \Mux36~2_combout ;
wire \Mux36~3_combout ;
wire \storeregister[24][27]~q ;
wire \Mux36~4_combout ;
wire \Mux36~5_combout ;
wire \Mux36~6_combout ;
wire \Mux36~0_combout ;
wire \Mux36~1_combout ;
wire \Mux36~7_combout ;
wire \Mux36~8_combout ;
wire \storeregister[13][27]~q ;
wire \Mux36~17_combout ;
wire \Mux36~18_combout ;
wire \Mux36~10_combout ;
wire \Mux36~11_combout ;
wire \Mux36~15_combout ;
wire \Mux36~12_combout ;
wire \storeregister[9][27]~feeder_combout ;
wire \storeregister[9][27]~q ;
wire \Mux36~13_combout ;
wire \Mux36~16_combout ;
wire \Mux45~7_combout ;
wire \Mux45~8_combout ;
wire \Mux45~0_combout ;
wire \Mux45~1_combout ;
wire \storeregister[26][18]~q ;
wire \Mux45~3_combout ;
wire \storeregister[16][18]~q ;
wire \Mux45~4_combout ;
wire \Mux45~5_combout ;
wire \Mux45~6_combout ;
wire \Mux45~12_combout ;
wire \Mux45~13_combout ;
wire \Mux45~15_combout ;
wire \Mux45~16_combout ;
wire \Mux45~10_combout ;
wire \Mux45~11_combout ;
wire \Mux45~17_combout ;
wire \Mux45~18_combout ;
wire \Mux46~7_combout ;
wire \Mux46~8_combout ;
wire \Mux46~0_combout ;
wire \Mux46~1_combout ;
wire \storeregister[22][17]~q ;
wire \Mux46~3_combout ;
wire \storeregister[28][17]~feeder_combout ;
wire \storeregister[28][17]~q ;
wire \Mux46~4_combout ;
wire \Mux46~5_combout ;
wire \Mux46~6_combout ;
wire \Mux46~17_combout ;
wire \Mux46~18_combout ;
wire \Mux46~14_combout ;
wire \Mux46~15_combout ;
wire \Mux46~12_combout ;
wire \Mux46~13_combout ;
wire \Mux46~16_combout ;
wire \Mux46~10_combout ;
wire \storeregister[9][17]~q ;
wire \Mux46~11_combout ;
wire \Mux47~0_combout ;
wire \Mux47~1_combout ;
wire \storeregister[19][16]~q ;
wire \Mux47~7_combout ;
wire \Mux47~8_combout ;
wire \storeregister[28][16]~feeder_combout ;
wire \storeregister[28][16]~q ;
wire \Mux47~5_combout ;
wire \Mux47~2_combout ;
wire \Mux47~3_combout ;
wire \Mux47~6_combout ;
wire \Mux47~12_combout ;
wire \Mux47~13_combout ;
wire \Mux47~14_combout ;
wire \storeregister[2][16]~q ;
wire \Mux47~15_combout ;
wire \Mux47~16_combout ;
wire \Mux47~10_combout ;
wire \storeregister[6][16]~q ;
wire \Mux47~11_combout ;
wire \Mux47~17_combout ;
wire \Mux47~18_combout ;
wire \storeregister[17][31]~q ;
wire \Mux32~0_combout ;
wire \Mux32~1_combout ;
wire \Mux32~7_combout ;
wire \Mux32~8_combout ;
wire \storeregister[16][31]~feeder_combout ;
wire \storeregister[16][31]~q ;
wire \Mux32~4_combout ;
wire \storeregister[28][31]~feeder_combout ;
wire \storeregister[28][31]~q ;
wire \Mux32~5_combout ;
wire \storeregister[22][31]~feeder_combout ;
wire \storeregister[22][31]~q ;
wire \Mux32~3_combout ;
wire \Mux32~6_combout ;
wire \storeregister[10][31]~q ;
wire \Mux32~10_combout ;
wire \Mux32~11_combout ;
wire \storeregister[13][31]~feeder_combout ;
wire \storeregister[13][31]~q ;
wire \Mux32~17_combout ;
wire \Mux32~18_combout ;
wire \Mux32~12_combout ;
wire \Mux32~13_combout ;
wire \Mux32~15_combout ;
wire \Mux32~16_combout ;
wire \Mux33~0_combout ;
wire \Mux33~1_combout ;
wire \Mux33~4_combout ;
wire \Mux33~5_combout ;
wire \storeregister[18][30]~q ;
wire \storeregister[22][30]~feeder_combout ;
wire \storeregister[22][30]~q ;
wire \Mux33~2_combout ;
wire \Mux33~3_combout ;
wire \Mux33~6_combout ;
wire \Mux33~7_combout ;
wire \Mux33~8_combout ;
wire \storeregister[5][30]~q ;
wire \Mux33~10_combout ;
wire \Mux33~11_combout ;
wire \Mux33~17_combout ;
wire \Mux33~18_combout ;
wire \storeregister[8][30]~q ;
wire \Mux33~12_combout ;
wire \Mux33~13_combout ;
wire \Mux33~14_combout ;
wire \Mux33~15_combout ;
wire \Mux33~16_combout ;
wire \Mux34~7_combout ;
wire \Mux34~8_combout ;
wire \Mux34~3_combout ;
wire \storeregister[28][29]~feeder_combout ;
wire \storeregister[28][29]~q ;
wire \storeregister[20][29]~feeder_combout ;
wire \storeregister[20][29]~q ;
wire \Mux34~5_combout ;
wire \Mux34~6_combout ;
wire \Mux34~0_combout ;
wire \Mux34~1_combout ;
wire \Mux34~10_combout ;
wire \Mux34~11_combout ;
wire \Mux34~13_combout ;
wire \storeregister[3][29]~q ;
wire \storeregister[1][29]~q ;
wire \Mux34~14_combout ;
wire \Mux34~15_combout ;
wire \Mux34~16_combout ;
wire \Mux34~17_combout ;
wire \Mux34~18_combout ;
wire \Mux35~7_combout ;
wire \Mux35~8_combout ;
wire \storeregister[18][28]~q ;
wire \storeregister[22][28]~feeder_combout ;
wire \storeregister[22][28]~q ;
wire \Mux35~2_combout ;
wire \Mux35~3_combout ;
wire \Mux35~4_combout ;
wire \Mux35~5_combout ;
wire \Mux35~6_combout ;
wire \Mux35~0_combout ;
wire \Mux35~1_combout ;
wire \storeregister[5][28]~q ;
wire \Mux35~10_combout ;
wire \Mux35~11_combout ;
wire \storeregister[1][28]~q ;
wire \Mux35~14_combout ;
wire \Mux35~15_combout ;
wire \Mux35~13_combout ;
wire \Mux35~16_combout ;
wire \Mux35~17_combout ;
wire \Mux35~18_combout ;
wire \storeregister[17][26]~q ;
wire \Mux37~0_combout ;
wire \Mux37~1_combout ;
wire \storeregister[18][26]~q ;
wire \Mux37~2_combout ;
wire \Mux37~3_combout ;
wire \storeregister[20][26]~q ;
wire \Mux37~4_combout ;
wire \Mux37~5_combout ;
wire \Mux37~6_combout ;
wire \Mux37~7_combout ;
wire \Mux37~8_combout ;
wire \storeregister[1][26]~q ;
wire \Mux37~14_combout ;
wire \Mux37~15_combout ;
wire \storeregister[8][26]~q ;
wire \Mux37~12_combout ;
wire \Mux37~13_combout ;
wire \Mux37~16_combout ;
wire \storeregister[5][26]~q ;
wire \storeregister[4][26]~q ;
wire \Mux37~10_combout ;
wire \Mux37~11_combout ;
wire \Mux37~17_combout ;
wire \Mux37~18_combout ;
wire \Mux38~7_combout ;
wire \Mux38~8_combout ;
wire \Mux38~0_combout ;
wire \Mux38~1_combout ;
wire \Mux38~3_combout ;
wire \storeregister[24][25]~q ;
wire \Mux38~4_combout ;
wire \Mux38~5_combout ;
wire \Mux38~6_combout ;
wire \Mux38~13_combout ;
wire \storeregister[1][25]~q ;
wire \Mux38~14_combout ;
wire \Mux38~15_combout ;
wire \Mux38~16_combout ;
wire \Mux38~17_combout ;
wire \Mux38~18_combout ;
wire \storeregister[10][25]~q ;
wire \Mux38~10_combout ;
wire \Mux38~11_combout ;
wire \storeregister[20][24]~feeder_combout ;
wire \storeregister[20][24]~q ;
wire \Mux39~4_combout ;
wire \Mux39~5_combout ;
wire \Mux39~3_combout ;
wire \Mux39~6_combout ;
wire \storeregister[17][24]~q ;
wire \Mux39~0_combout ;
wire \Mux39~1_combout ;
wire \storeregister[23][24]~feeder_combout ;
wire \storeregister[23][24]~q ;
wire \Mux39~7_combout ;
wire \Mux39~8_combout ;
wire \storeregister[5][24]~q ;
wire \Mux39~10_combout ;
wire \storeregister[6][24]~q ;
wire \Mux39~11_combout ;
wire \storeregister[12][24]~q ;
wire \Mux39~17_combout ;
wire \Mux39~18_combout ;
wire \Mux39~12_combout ;
wire \Mux39~13_combout ;
wire \storeregister[1][24]~q ;
wire \Mux39~14_combout ;
wire \Mux39~15_combout ;
wire \Mux39~16_combout ;
wire \Mux40~4_combout ;
wire \Mux40~5_combout ;
wire \storeregister[22][23]~q ;
wire \storeregister[18][23]~q ;
wire \Mux40~2_combout ;
wire \Mux40~3_combout ;
wire \Mux40~6_combout ;
wire \Mux40~7_combout ;
wire \Mux40~8_combout ;
wire \Mux40~0_combout ;
wire \Mux40~1_combout ;
wire \Mux40~17_combout ;
wire \Mux40~18_combout ;
wire \Mux40~13_combout ;
wire \Mux40~14_combout ;
wire \Mux40~15_combout ;
wire \Mux40~16_combout ;
wire \storeregister[8][23]~q ;
wire \storeregister[10][23]~q ;
wire \Mux40~10_combout ;
wire \Mux40~11_combout ;
wire \Mux41~7_combout ;
wire \Mux41~8_combout ;
wire \storeregister[20][22]~q ;
wire \Mux41~4_combout ;
wire \Mux41~5_combout ;
wire \Mux41~2_combout ;
wire \Mux41~3_combout ;
wire \Mux41~6_combout ;
wire \storeregister[21][22]~feeder_combout ;
wire \storeregister[21][22]~q ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \Mux41~17_combout ;
wire \Mux41~18_combout ;
wire \Mux41~10_combout ;
wire \Mux41~11_combout ;
wire \storeregister[8][22]~q ;
wire \Mux41~12_combout ;
wire \Mux41~13_combout ;
wire \storeregister[3][22]~q ;
wire \storeregister[1][22]~q ;
wire \Mux41~14_combout ;
wire \Mux41~15_combout ;
wire \Mux41~16_combout ;
wire \Mux42~7_combout ;
wire \Mux42~8_combout ;
wire \storeregister[20][21]~q ;
wire \storeregister[16][21]~q ;
wire \Mux42~4_combout ;
wire \Mux42~5_combout ;
wire \storeregister[30][21]~q ;
wire \Mux42~3_combout ;
wire \Mux42~6_combout ;
wire \Mux42~0_combout ;
wire \Mux42~1_combout ;
wire \Mux42~14_combout ;
wire \storeregister[2][21]~q ;
wire \Mux42~15_combout ;
wire \Mux42~12_combout ;
wire \Mux42~13_combout ;
wire \Mux42~16_combout ;
wire \Mux42~17_combout ;
wire \Mux42~18_combout ;
wire \storeregister[9][21]~q ;
wire \Mux42~10_combout ;
wire \Mux42~11_combout ;
wire \Mux43~0_combout ;
wire \Mux43~1_combout ;
wire \Mux43~3_combout ;
wire \Mux43~4_combout ;
wire \storeregister[24][20]~q ;
wire \Mux43~5_combout ;
wire \Mux43~6_combout ;
wire \storeregister[23][20]~feeder_combout ;
wire \storeregister[23][20]~q ;
wire \Mux43~7_combout ;
wire \Mux43~8_combout ;
wire \Mux43~10_combout ;
wire \Mux43~11_combout ;
wire \storeregister[1][20]~q ;
wire \storeregister[3][20]~q ;
wire \Mux43~14_combout ;
wire \Mux43~15_combout ;
wire \Mux43~12_combout ;
wire \Mux43~13_combout ;
wire \Mux43~16_combout ;
wire \Mux43~17_combout ;
wire \Mux43~18_combout ;
wire \Mux44~7_combout ;
wire \Mux44~8_combout ;
wire \Mux44~0_combout ;
wire \Mux44~1_combout ;
wire \storeregister[26][19]~feeder_combout ;
wire \storeregister[26][19]~q ;
wire \Mux44~2_combout ;
wire \Mux44~3_combout ;
wire \storeregister[24][19]~feeder_combout ;
wire \storeregister[24][19]~q ;
wire \Mux44~4_combout ;
wire \Mux44~5_combout ;
wire \Mux44~6_combout ;
wire \storeregister[10][19]~q ;
wire \Mux44~10_combout ;
wire \Mux44~11_combout ;
wire \Mux44~14_combout ;
wire \Mux44~15_combout ;
wire \storeregister[4][19]~q ;
wire \Mux44~12_combout ;
wire \Mux44~13_combout ;
wire \Mux44~16_combout ;
wire \Mux44~17_combout ;
wire \Mux44~18_combout ;
wire \storeregister[18][10]~q ;
wire \Mux53~2_combout ;
wire \Mux53~3_combout ;
wire \storeregister[16][10]~q ;
wire \storeregister[24][10]~q ;
wire \Mux53~4_combout ;
wire \Mux53~5_combout ;
wire \Mux53~6_combout ;
wire \Mux53~7_combout ;
wire \Mux53~8_combout ;
wire \Mux53~0_combout ;
wire \Mux53~1_combout ;
wire \Mux53~17_combout ;
wire \Mux53~18_combout ;
wire \Mux53~10_combout ;
wire \Mux53~11_combout ;
wire \storeregister[6][10]~q ;
wire \Mux53~12_combout ;
wire \Mux53~13_combout ;
wire \storeregister[1][10]~q ;
wire \Mux53~14_combout ;
wire \Mux53~15_combout ;
wire \Mux53~16_combout ;
wire \Mux49~7_combout ;
wire \Mux49~8_combout ;
wire \Mux49~0_combout ;
wire \Mux49~1_combout ;
wire \Mux49~2_combout ;
wire \Mux49~3_combout ;
wire \Mux49~5_combout ;
wire \Mux49~6_combout ;
wire \Mux49~17_combout ;
wire \Mux49~18_combout ;
wire \Mux49~12_combout ;
wire \Mux49~13_combout ;
wire \storeregister[3][14]~q ;
wire \storeregister[1][14]~q ;
wire \Mux49~14_combout ;
wire \Mux49~15_combout ;
wire \Mux49~16_combout ;
wire \storeregister[5][14]~q ;
wire \storeregister[4][14]~q ;
wire \Mux49~10_combout ;
wire \Mux49~11_combout ;
wire \Mux54~7_combout ;
wire \Mux54~8_combout ;
wire \Mux54~0_combout ;
wire \storeregister[25][9]~feeder_combout ;
wire \storeregister[25][9]~q ;
wire \Mux54~1_combout ;
wire \storeregister[22][9]~q ;
wire \Mux54~3_combout ;
wire \storeregister[16][9]~q ;
wire \Mux54~4_combout ;
wire \storeregister[20][9]~feeder_combout ;
wire \storeregister[20][9]~q ;
wire \Mux54~5_combout ;
wire \Mux54~6_combout ;
wire \Mux54~17_combout ;
wire \Mux54~18_combout ;
wire \storeregister[4][9]~q ;
wire \Mux54~12_combout ;
wire \Mux54~13_combout ;
wire \storeregister[1][9]~q ;
wire \Mux54~14_combout ;
wire \Mux54~15_combout ;
wire \Mux54~16_combout ;
wire \Mux54~10_combout ;
wire \Mux54~11_combout ;
wire \Mux55~7_combout ;
wire \Mux55~8_combout ;
wire \Mux55~0_combout ;
wire \Mux55~1_combout ;
wire \storeregister[22][8]~q ;
wire \Mux55~2_combout ;
wire \Mux55~3_combout ;
wire \storeregister[24][8]~feeder_combout ;
wire \storeregister[24][8]~q ;
wire \Mux55~5_combout ;
wire \Mux55~6_combout ;
wire \Mux55~17_combout ;
wire \Mux55~18_combout ;
wire \storeregister[5][8]~q ;
wire \storeregister[4][8]~q ;
wire \Mux55~10_combout ;
wire \Mux55~11_combout ;
wire \Mux55~12_combout ;
wire \Mux55~13_combout ;
wire \storeregister[3][8]~q ;
wire \storeregister[1][8]~q ;
wire \Mux55~14_combout ;
wire \Mux55~15_combout ;
wire \Mux55~16_combout ;
wire \Mux56~0_combout ;
wire \Mux56~1_combout ;
wire \Mux56~7_combout ;
wire \Mux56~8_combout ;
wire \Mux56~4_combout ;
wire \Mux56~5_combout ;
wire \Mux56~3_combout ;
wire \Mux56~6_combout ;
wire \Mux56~17_combout ;
wire \Mux56~18_combout ;
wire \Mux56~14_combout ;
wire \Mux56~15_combout ;
wire \Mux56~13_combout ;
wire \Mux56~16_combout ;
wire \storeregister[11][7]~feeder_combout ;
wire \storeregister[11][7]~q ;
wire \Mux56~10_combout ;
wire \Mux56~11_combout ;
wire \Mux57~7_combout ;
wire \Mux57~8_combout ;
wire \Mux57~2_combout ;
wire \Mux57~3_combout ;
wire \Mux57~5_combout ;
wire \Mux57~6_combout ;
wire \storeregister[17][6]~q ;
wire \Mux57~0_combout ;
wire \Mux57~1_combout ;
wire \Mux57~12_combout ;
wire \Mux57~13_combout ;
wire \Mux57~14_combout ;
wire \Mux57~15_combout ;
wire \Mux57~16_combout ;
wire \storeregister[4][6]~q ;
wire \storeregister[5][6]~q ;
wire \Mux57~10_combout ;
wire \Mux57~11_combout ;
wire \Mux57~17_combout ;
wire \Mux57~18_combout ;
wire \Mux58~0_combout ;
wire \Mux58~1_combout ;
wire \Mux58~7_combout ;
wire \Mux58~8_combout ;
wire \storeregister[16][5]~q ;
wire \storeregister[24][5]~feeder_combout ;
wire \storeregister[24][5]~q ;
wire \Mux58~4_combout ;
wire \Mux58~5_combout ;
wire \storeregister[22][5]~feeder_combout ;
wire \storeregister[22][5]~q ;
wire \storeregister[30][5]~q ;
wire \Mux58~3_combout ;
wire \Mux58~6_combout ;
wire \Mux58~17_combout ;
wire \Mux58~18_combout ;
wire \storeregister[10][5]~q ;
wire \Mux58~10_combout ;
wire \Mux58~11_combout ;
wire \Mux58~12_combout ;
wire \Mux58~13_combout ;
wire \Mux58~14_combout ;
wire \Mux58~15_combout ;
wire \Mux58~16_combout ;
wire \Mux50~7_combout ;
wire \Mux50~8_combout ;
wire \Mux50~3_combout ;
wire \storeregister[16][13]~feeder_combout ;
wire \storeregister[16][13]~q ;
wire \Mux50~4_combout ;
wire \Mux50~5_combout ;
wire \Mux50~6_combout ;
wire \storeregister[17][13]~q ;
wire \Mux50~0_combout ;
wire \Mux50~1_combout ;
wire \storeregister[10][13]~q ;
wire \Mux50~10_combout ;
wire \Mux50~11_combout ;
wire \Mux50~14_combout ;
wire \Mux50~15_combout ;
wire \storeregister[4][13]~q ;
wire \Mux50~12_combout ;
wire \Mux50~13_combout ;
wire \Mux50~16_combout ;
wire \Mux50~17_combout ;
wire \Mux50~18_combout ;
wire \storeregister[27][11]~feeder_combout ;
wire \storeregister[27][11]~q ;
wire \Mux52~7_combout ;
wire \Mux52~8_combout ;
wire \Mux52~2_combout ;
wire \Mux52~3_combout ;
wire \storeregister[24][11]~q ;
wire \Mux52~4_combout ;
wire \storeregister[20][11]~feeder_combout ;
wire \storeregister[20][11]~q ;
wire \Mux52~5_combout ;
wire \Mux52~6_combout ;
wire \Mux52~0_combout ;
wire \Mux52~1_combout ;
wire \Mux52~12_combout ;
wire \Mux52~13_combout ;
wire \Mux52~15_combout ;
wire \Mux52~16_combout ;
wire \Mux52~17_combout ;
wire \Mux52~18_combout ;
wire \storeregister[10][11]~q ;
wire \Mux52~10_combout ;
wire \Mux52~11_combout ;


// Location: FF_X49_Y36_N3
dffeas \storeregister[22][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][1] .is_wysiwyg = "true";
defparam \storeregister[22][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N9
dffeas \storeregister[18][1] (
	.clk(!CLK),
	.d(\storeregister[18][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][1] .is_wysiwyg = "true";
defparam \storeregister[18][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N2
cycloneive_lcell_comb \Mux62~2 (
// Equation(s):
// \Mux62~2_combout  = (temp_imemload_output_18 & ((\storeregister[22][1]~q ) # ((temp_imemload_output_19)))) # (!temp_imemload_output_18 & (((\storeregister[18][1]~q  & !temp_imemload_output_19))))

	.dataa(\storeregister[22][1]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[18][1]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux62~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~2 .lut_mask = 16'hCCB8;
defparam \Mux62~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N18
cycloneive_lcell_comb \Mux62~12 (
// Equation(s):
// \Mux62~12_combout  = (temp_imemload_output_16 & (temp_imemload_output_17)) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[10][1]~q ))) # (!temp_imemload_output_17 & (\storeregister[8][1]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[8][1]~q ),
	.datad(\storeregister[10][1]~q ),
	.cin(gnd),
	.combout(\Mux62~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~12 .lut_mask = 16'hDC98;
defparam \Mux62~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N2
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (temp_imemload_output_23 & (((\storeregister[22][1]~q ) # (temp_imemload_output_24)))) # (!temp_imemload_output_23 & (\storeregister[18][1]~q  & ((!temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[18][1]~q ),
	.datac(\storeregister[22][1]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'hAAE4;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N2
cycloneive_lcell_comb \Mux30~4 (
// Equation(s):
// \Mux30~4_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\storeregister[20][1]~q )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & (\storeregister[16][1]~q )))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][1]~q ),
	.datad(\storeregister[20][1]~q ),
	.cin(gnd),
	.combout(\Mux30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~4 .lut_mask = 16'hBA98;
defparam \Mux30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N12
cycloneive_lcell_comb \Mux30~14 (
// Equation(s):
// \Mux30~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][1]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][1]~q ))))

	.dataa(\storeregister[1][1]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[3][1]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux30~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~14 .lut_mask = 16'hE200;
defparam \Mux30~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N25
dffeas \storeregister[26][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][0] .is_wysiwyg = "true";
defparam \storeregister[26][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N3
dffeas \storeregister[18][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][0] .is_wysiwyg = "true";
defparam \storeregister[18][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N24
cycloneive_lcell_comb \Mux63~2 (
// Equation(s):
// \Mux63~2_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\storeregister[26][0]~q )) # (!temp_imemload_output_19 & ((\storeregister[18][0]~q )))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[26][0]~q ),
	.datad(\storeregister[18][0]~q ),
	.cin(gnd),
	.combout(\Mux63~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~2 .lut_mask = 16'hD9C8;
defparam \Mux63~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N30
cycloneive_lcell_comb \Mux63~4 (
// Equation(s):
// \Mux63~4_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\storeregister[24][0]~q )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & (\storeregister[16][0]~q )))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[16][0]~q ),
	.datad(\storeregister[24][0]~q ),
	.cin(gnd),
	.combout(\Mux63~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~4 .lut_mask = 16'hBA98;
defparam \Mux63~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N16
cycloneive_lcell_comb \Mux63~12 (
// Equation(s):
// \Mux63~12_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[5][0]~q ))) # (!temp_imemload_output_16 & (\storeregister[4][0]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[4][0]~q ),
	.datac(\storeregister[5][0]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux63~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~12 .lut_mask = 16'hFA44;
defparam \Mux63~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N7
dffeas \storeregister[1][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][0] .is_wysiwyg = "true";
defparam \storeregister[1][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N6
cycloneive_lcell_comb \Mux63~14 (
// Equation(s):
// \Mux63~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[3][0]~q ))) # (!temp_imemload_output_17 & (\storeregister[1][0]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[1][0]~q ),
	.datad(\storeregister[3][0]~q ),
	.cin(gnd),
	.combout(\Mux63~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~14 .lut_mask = 16'hA820;
defparam \Mux63~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N2
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (temp_imemload_output_24 & ((\storeregister[26][0]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[18][0]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[26][0]~q ),
	.datac(\storeregister[18][0]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hAAD8;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N7
dffeas \storeregister[28][2] (
	.clk(!CLK),
	.d(\storeregister[28][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][2] .is_wysiwyg = "true";
defparam \storeregister[28][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N13
dffeas \storeregister[30][3] (
	.clk(!CLK),
	.d(\storeregister[30][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][3] .is_wysiwyg = "true";
defparam \storeregister[30][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N14
cycloneive_lcell_comb \Mux28~14 (
// Equation(s):
// \Mux28~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][3]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][3]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[1][3]~q ),
	.datad(\storeregister[3][3]~q ),
	.cin(gnd),
	.combout(\Mux28~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~14 .lut_mask = 16'hA820;
defparam \Mux28~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N21
dffeas \storeregister[16][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][8] .is_wysiwyg = "true";
defparam \storeregister[16][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N14
cycloneive_lcell_comb \Mux23~4 (
// Equation(s):
// \Mux23~4_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23) # (\storeregister[24][8]~q )))) # (!temp_imemload_output_24 & (\storeregister[16][8]~q  & (!temp_imemload_output_23)))

	.dataa(\storeregister[16][8]~q ),
	.datab(temp_imemload_output_24),
	.datac(temp_imemload_output_23),
	.datad(\storeregister[24][8]~q ),
	.cin(gnd),
	.combout(\Mux23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~4 .lut_mask = 16'hCEC2;
defparam \Mux23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N10
cycloneive_lcell_comb \Mux23~12 (
// Equation(s):
// \Mux23~12_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[5][8]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[4][8]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[4][8]~q ),
	.datad(\storeregister[5][8]~q ),
	.cin(gnd),
	.combout(\Mux23~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~12 .lut_mask = 16'hBA98;
defparam \Mux23~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N2
cycloneive_lcell_comb \Mux23~14 (
// Equation(s):
// \Mux23~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][8]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][8]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[1][8]~q ),
	.datad(\storeregister[3][8]~q ),
	.cin(gnd),
	.combout(\Mux23~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~14 .lut_mask = 16'hA820;
defparam \Mux23~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N5
dffeas \storeregister[26][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][7] .is_wysiwyg = "true";
defparam \storeregister[26][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N14
cycloneive_lcell_comb \Mux25~12 (
// Equation(s):
// \Mux25~12_combout  = (temp_imemload_output_21 & ((\storeregister[5][6]~q ) # ((temp_imemload_output_22)))) # (!temp_imemload_output_21 & (((\storeregister[4][6]~q  & !temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[5][6]~q ),
	.datac(\storeregister[4][6]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux25~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~12 .lut_mask = 16'hAAD8;
defparam \Mux25~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N27
dffeas \storeregister[8][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][5] .is_wysiwyg = "true";
defparam \storeregister[8][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N26
cycloneive_lcell_comb \Mux26~12 (
// Equation(s):
// \Mux26~12_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\storeregister[10][5]~q )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & (\storeregister[8][5]~q )))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[8][5]~q ),
	.datad(\storeregister[10][5]~q ),
	.cin(gnd),
	.combout(\Mux26~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~12 .lut_mask = 16'hBA98;
defparam \Mux26~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N18
cycloneive_lcell_comb \Mux17~12 (
// Equation(s):
// \Mux17~12_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[5][14]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[4][14]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[4][14]~q ),
	.datad(\storeregister[5][14]~q ),
	.cin(gnd),
	.combout(\Mux17~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~12 .lut_mask = 16'hBA98;
defparam \Mux17~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N6
cycloneive_lcell_comb \Mux17~14 (
// Equation(s):
// \Mux17~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[3][14]~q )) # (!temp_imemload_output_22 & ((\storeregister[1][14]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[3][14]~q ),
	.datac(\storeregister[1][14]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux17~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~14 .lut_mask = 16'h88A0;
defparam \Mux17~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N8
cycloneive_lcell_comb \Mux16~4 (
// Equation(s):
// \Mux16~4_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\storeregister[20][15]~q )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & ((\storeregister[16][15]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[20][15]~q ),
	.datad(\storeregister[16][15]~q ),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~4 .lut_mask = 16'hB9A8;
defparam \Mux16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N16
cycloneive_lcell_comb \Mux16~12 (
// Equation(s):
// \Mux16~12_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22)))) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[10][15]~q )) # (!temp_imemload_output_22 & ((\storeregister[8][15]~q )))))

	.dataa(\storeregister[10][15]~q ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[8][15]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux16~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~12 .lut_mask = 16'hEE30;
defparam \Mux16~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N13
dffeas \storeregister[20][13] (
	.clk(!CLK),
	.d(\storeregister[20][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][13] .is_wysiwyg = "true";
defparam \storeregister[20][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N10
cycloneive_lcell_comb \Mux18~4 (
// Equation(s):
// \Mux18~4_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\storeregister[20][13]~q )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & (\storeregister[16][13]~q )))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][13]~q ),
	.datad(\storeregister[20][13]~q ),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~4 .lut_mask = 16'hBA98;
defparam \Mux18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N15
dffeas \storeregister[8][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][13] .is_wysiwyg = "true";
defparam \storeregister[8][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N14
cycloneive_lcell_comb \Mux18~12 (
// Equation(s):
// \Mux18~12_combout  = (temp_imemload_output_22 & ((\storeregister[10][13]~q ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((\storeregister[8][13]~q  & !temp_imemload_output_21))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[10][13]~q ),
	.datac(\storeregister[8][13]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux18~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~12 .lut_mask = 16'hAAD8;
defparam \Mux18~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N18
cycloneive_lcell_comb \Mux19~12 (
// Equation(s):
// \Mux19~12_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & (\storeregister[5][12]~q )) # (!temp_imemload_output_21 & ((\storeregister[4][12]~q )))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[5][12]~q ),
	.datac(\storeregister[4][12]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux19~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~12 .lut_mask = 16'hEE50;
defparam \Mux19~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N0
cycloneive_lcell_comb \Mux21~4 (
// Equation(s):
// \Mux21~4_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[24][10]~q )) # (!temp_imemload_output_24 & ((\storeregister[16][10]~q )))))

	.dataa(\storeregister[24][10]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[16][10]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~4 .lut_mask = 16'hEE30;
defparam \Mux21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N17
dffeas \storeregister[30][11] (
	.clk(!CLK),
	.d(\storeregister[30][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][11] .is_wysiwyg = "true";
defparam \storeregister[30][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N11
dffeas \storeregister[8][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][11] .is_wysiwyg = "true";
defparam \storeregister[8][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N10
cycloneive_lcell_comb \Mux20~12 (
// Equation(s):
// \Mux20~12_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\storeregister[10][11]~q )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & (\storeregister[8][11]~q )))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[8][11]~q ),
	.datad(\storeregister[10][11]~q ),
	.cin(gnd),
	.combout(\Mux20~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~12 .lut_mask = 16'hBA98;
defparam \Mux20~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N31
dffeas \storeregister[1][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][11] .is_wysiwyg = "true";
defparam \storeregister[1][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N15
dffeas \storeregister[18][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][9] .is_wysiwyg = "true";
defparam \storeregister[18][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N4
cycloneive_lcell_comb \Mux22~2 (
// Equation(s):
// \Mux22~2_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[22][9]~q )) # (!temp_imemload_output_23 & ((\storeregister[18][9]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[22][9]~q ),
	.datad(\storeregister[18][9]~q ),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~2 .lut_mask = 16'hD9C8;
defparam \Mux22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N10
cycloneive_lcell_comb \Mux22~4 (
// Equation(s):
// \Mux22~4_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24) # (\storeregister[20][9]~q )))) # (!temp_imemload_output_23 & (\storeregister[16][9]~q  & (!temp_imemload_output_24)))

	.dataa(\storeregister[16][9]~q ),
	.datab(temp_imemload_output_23),
	.datac(temp_imemload_output_24),
	.datad(\storeregister[20][9]~q ),
	.cin(gnd),
	.combout(\Mux22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~4 .lut_mask = 16'hCEC2;
defparam \Mux22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N10
cycloneive_lcell_comb \Mux59~2 (
// Equation(s):
// \Mux59~2_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[22][4]~q ))) # (!temp_imemload_output_18 & (\storeregister[18][4]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[18][4]~q ),
	.datad(\storeregister[22][4]~q ),
	.cin(gnd),
	.combout(\Mux59~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~2 .lut_mask = 16'hDC98;
defparam \Mux59~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N12
cycloneive_lcell_comb \Mux59~4 (
// Equation(s):
// \Mux59~4_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\storeregister[20][4]~q )) # (!temp_imemload_output_18 & ((\storeregister[16][4]~q )))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[20][4]~q ),
	.datad(\storeregister[16][4]~q ),
	.cin(gnd),
	.combout(\Mux59~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~4 .lut_mask = 16'hD9C8;
defparam \Mux59~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N14
cycloneive_lcell_comb \Mux59~12 (
// Equation(s):
// \Mux59~12_combout  = (temp_imemload_output_16 & (temp_imemload_output_17)) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[10][4]~q ))) # (!temp_imemload_output_17 & (\storeregister[8][4]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[8][4]~q ),
	.datad(\storeregister[10][4]~q ),
	.cin(gnd),
	.combout(\Mux59~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~12 .lut_mask = 16'hDC98;
defparam \Mux59~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N3
dffeas \storeregister[18][31] (
	.clk(!CLK),
	.d(\storeregister[18][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][31] .is_wysiwyg = "true";
defparam \storeregister[18][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N12
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[22][31]~q ))) # (!temp_imemload_output_23 & (\storeregister[18][31]~q ))))

	.dataa(\storeregister[18][31]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[22][31]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hFC22;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N11
dffeas \storeregister[8][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][31] .is_wysiwyg = "true";
defparam \storeregister[8][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N10
cycloneive_lcell_comb \Mux0~12 (
// Equation(s):
// \Mux0~12_combout  = (temp_imemload_output_22 & ((\storeregister[10][31]~q ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((\storeregister[8][31]~q  & !temp_imemload_output_21))))

	.dataa(\storeregister[10][31]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[8][31]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~12 .lut_mask = 16'hCCB8;
defparam \Mux0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N27
dffeas \storeregister[1][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][31] .is_wysiwyg = "true";
defparam \storeregister[1][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N31
dffeas \storeregister[4][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][30] .is_wysiwyg = "true";
defparam \storeregister[4][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N30
cycloneive_lcell_comb \Mux1~12 (
// Equation(s):
// \Mux1~12_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[5][30]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[4][30]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[4][30]~q ),
	.datad(\storeregister[5][30]~q ),
	.cin(gnd),
	.combout(\Mux1~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~12 .lut_mask = 16'hBA98;
defparam \Mux1~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N20
cycloneive_lcell_comb \Mux2~14 (
// Equation(s):
// \Mux2~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][29]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][29]~q ))))

	.dataa(\storeregister[1][29]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[3][29]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~14 .lut_mask = 16'hE200;
defparam \Mux2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N2
cycloneive_lcell_comb \Mux5~12 (
// Equation(s):
// \Mux5~12_combout  = (temp_imemload_output_21 & ((\storeregister[5][26]~q ) # ((temp_imemload_output_22)))) # (!temp_imemload_output_21 & (((\storeregister[4][26]~q  & !temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[5][26]~q ),
	.datac(\storeregister[4][26]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux5~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~12 .lut_mask = 16'hAAD8;
defparam \Mux5~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N1
dffeas \storeregister[26][25] (
	.clk(!CLK),
	.d(\storeregister[26][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][25] .is_wysiwyg = "true";
defparam \storeregister[26][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y41_N31
dffeas \storeregister[4][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][25] .is_wysiwyg = "true";
defparam \storeregister[4][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y39_N13
dffeas \storeregister[8][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][25] .is_wysiwyg = "true";
defparam \storeregister[8][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N12
cycloneive_lcell_comb \Mux6~12 (
// Equation(s):
// \Mux6~12_combout  = (temp_imemload_output_22 & ((\storeregister[10][25]~q ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((\storeregister[8][25]~q  & !temp_imemload_output_21))))

	.dataa(\storeregister[10][25]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[8][25]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux6~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~12 .lut_mask = 16'hCCB8;
defparam \Mux6~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N13
dffeas \storeregister[28][28] (
	.clk(!CLK),
	.d(\storeregister[28][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][28] .is_wysiwyg = "true";
defparam \storeregister[28][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N31
dffeas \storeregister[8][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][28] .is_wysiwyg = "true";
defparam \storeregister[8][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y41_N27
dffeas \storeregister[4][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][28] .is_wysiwyg = "true";
defparam \storeregister[4][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N26
cycloneive_lcell_comb \Mux3~12 (
// Equation(s):
// \Mux3~12_combout  = (temp_imemload_output_22 & (temp_imemload_output_21)) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[5][28]~q ))) # (!temp_imemload_output_21 & (\storeregister[4][28]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[4][28]~q ),
	.datad(\storeregister[5][28]~q ),
	.cin(gnd),
	.combout(\Mux3~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~12 .lut_mask = 16'hDC98;
defparam \Mux3~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N12
cycloneive_lcell_comb \Mux4~2 (
// Equation(s):
// \Mux4~2_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[22][27]~q )) # (!temp_imemload_output_23 & ((\storeregister[18][27]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[22][27]~q ),
	.datad(\storeregister[18][27]~q ),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~2 .lut_mask = 16'hD9C8;
defparam \Mux4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N13
dffeas \storeregister[18][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][17] .is_wysiwyg = "true";
defparam \storeregister[18][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N22
cycloneive_lcell_comb \Mux14~2 (
// Equation(s):
// \Mux14~2_combout  = (temp_imemload_output_23 & (((\storeregister[22][17]~q ) # (temp_imemload_output_24)))) # (!temp_imemload_output_23 & (\storeregister[18][17]~q  & ((!temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[18][17]~q ),
	.datac(\storeregister[22][17]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~2 .lut_mask = 16'hAAE4;
defparam \Mux14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N23
dffeas \storeregister[20][17] (
	.clk(!CLK),
	.d(\storeregister[20][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][17] .is_wysiwyg = "true";
defparam \storeregister[20][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N27
dffeas \storeregister[16][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][20] .is_wysiwyg = "true";
defparam \storeregister[16][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N26
cycloneive_lcell_comb \Mux11~4 (
// Equation(s):
// \Mux11~4_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[24][20]~q ))) # (!temp_imemload_output_24 & (\storeregister[16][20]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][20]~q ),
	.datad(\storeregister[24][20]~q ),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~4 .lut_mask = 16'hDC98;
defparam \Mux11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N28
cycloneive_lcell_comb \Mux11~14 (
// Equation(s):
// \Mux11~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][20]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][20]~q ))))

	.dataa(\storeregister[1][20]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[3][20]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux11~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~14 .lut_mask = 16'hE200;
defparam \Mux11~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N31
dffeas \storeregister[8][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][19] .is_wysiwyg = "true";
defparam \storeregister[8][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N30
cycloneive_lcell_comb \Mux12~12 (
// Equation(s):
// \Mux12~12_combout  = (temp_imemload_output_22 & ((\storeregister[10][19]~q ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((\storeregister[8][19]~q  & !temp_imemload_output_21))))

	.dataa(\storeregister[10][19]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[8][19]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux12~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~12 .lut_mask = 16'hCCB8;
defparam \Mux12~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N27
dffeas \storeregister[18][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][18] .is_wysiwyg = "true";
defparam \storeregister[18][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N26
cycloneive_lcell_comb \Mux13~2 (
// Equation(s):
// \Mux13~2_combout  = (temp_imemload_output_24 & ((\storeregister[26][18]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[18][18]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[26][18]~q ),
	.datac(\storeregister[18][18]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~2 .lut_mask = 16'hAAD8;
defparam \Mux13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N13
dffeas \storeregister[3][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][18] .is_wysiwyg = "true";
defparam \storeregister[3][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N3
dffeas \storeregister[1][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][18] .is_wysiwyg = "true";
defparam \storeregister[1][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N12
cycloneive_lcell_comb \Mux13~14 (
// Equation(s):
// \Mux13~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][18]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][18]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[1][18]~q ),
	.datac(\storeregister[3][18]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux13~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~14 .lut_mask = 16'hE400;
defparam \Mux13~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N21
dffeas \storeregister[22][24] (
	.clk(!CLK),
	.d(\storeregister[22][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][24] .is_wysiwyg = "true";
defparam \storeregister[22][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N2
cycloneive_lcell_comb \Mux8~2 (
// Equation(s):
// \Mux8~2_combout  = (temp_imemload_output_23 & ((\storeregister[22][23]~q ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\storeregister[18][23]~q  & !temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[22][23]~q ),
	.datac(\storeregister[18][23]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~2 .lut_mask = 16'hAAD8;
defparam \Mux8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N8
cycloneive_lcell_comb \Mux8~12 (
// Equation(s):
// \Mux8~12_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[10][23]~q ))) # (!temp_imemload_output_22 & (\storeregister[8][23]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[8][23]~q ),
	.datad(\storeregister[10][23]~q ),
	.cin(gnd),
	.combout(\Mux8~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~12 .lut_mask = 16'hDC98;
defparam \Mux8~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N21
dffeas \storeregister[26][22] (
	.clk(!CLK),
	.d(\storeregister[26][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][22] .is_wysiwyg = "true";
defparam \storeregister[26][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N3
dffeas \storeregister[18][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][22] .is_wysiwyg = "true";
defparam \storeregister[18][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N2
cycloneive_lcell_comb \Mux9~2 (
// Equation(s):
// \Mux9~2_combout  = (temp_imemload_output_24 & ((\storeregister[26][22]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[18][22]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[26][22]~q ),
	.datac(\storeregister[18][22]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~2 .lut_mask = 16'hAAD8;
defparam \Mux9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N16
cycloneive_lcell_comb \Mux9~14 (
// Equation(s):
// \Mux9~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][22]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][22]~q ))))

	.dataa(\storeregister[1][22]~q ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[3][22]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux9~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~14 .lut_mask = 16'hC088;
defparam \Mux9~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N30
cycloneive_lcell_comb \Mux10~4 (
// Equation(s):
// \Mux10~4_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\storeregister[20][21]~q )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & ((\storeregister[16][21]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[20][21]~q ),
	.datad(\storeregister[16][21]~q ),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~4 .lut_mask = 16'hB9A8;
defparam \Mux10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N14
cycloneive_lcell_comb \Mux48~2 (
// Equation(s):
// \Mux48~2_combout  = (temp_imemload_output_19 & ((\storeregister[26][15]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\storeregister[18][15]~q  & !temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[26][15]~q ),
	.datac(\storeregister[18][15]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux48~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~2 .lut_mask = 16'hAAD8;
defparam \Mux48~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N10
cycloneive_lcell_comb \Mux36~14 (
// Equation(s):
// \Mux36~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][27]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][27]~q )))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[3][27]~q ),
	.datac(\storeregister[1][27]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux36~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~14 .lut_mask = 16'h88A0;
defparam \Mux36~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N22
cycloneive_lcell_comb \Mux45~2 (
// Equation(s):
// \Mux45~2_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\storeregister[22][18]~q )) # (!temp_imemload_output_18 & ((\storeregister[18][18]~q )))))

	.dataa(\storeregister[22][18]~q ),
	.datab(\storeregister[18][18]~q ),
	.datac(temp_imemload_output_19),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux45~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~2 .lut_mask = 16'hFA0C;
defparam \Mux45~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N2
cycloneive_lcell_comb \Mux45~14 (
// Equation(s):
// \Mux45~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[3][18]~q ))) # (!temp_imemload_output_17 & (\storeregister[1][18]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[1][18]~q ),
	.datad(\storeregister[3][18]~q ),
	.cin(gnd),
	.combout(\Mux45~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~14 .lut_mask = 16'hA820;
defparam \Mux45~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N12
cycloneive_lcell_comb \Mux46~2 (
// Equation(s):
// \Mux46~2_combout  = (temp_imemload_output_19 & ((\storeregister[26][17]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\storeregister[18][17]~q  & !temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[26][17]~q ),
	.datac(\storeregister[18][17]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~2 .lut_mask = 16'hAAD8;
defparam \Mux46~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N12
cycloneive_lcell_comb \Mux47~4 (
// Equation(s):
// \Mux47~4_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[20][16]~q ))) # (!temp_imemload_output_18 & (\storeregister[16][16]~q ))))

	.dataa(\storeregister[16][16]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[20][16]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux47~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~4 .lut_mask = 16'hFC22;
defparam \Mux47~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N4
cycloneive_lcell_comb \Mux32~2 (
// Equation(s):
// \Mux32~2_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\storeregister[26][31]~q )) # (!temp_imemload_output_19 & ((\storeregister[18][31]~q )))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[26][31]~q ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[18][31]~q ),
	.cin(gnd),
	.combout(\Mux32~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~2 .lut_mask = 16'hE5E0;
defparam \Mux32~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N26
cycloneive_lcell_comb \Mux32~14 (
// Equation(s):
// \Mux32~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][31]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][31]~q )))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[3][31]~q ),
	.datac(\storeregister[1][31]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux32~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~14 .lut_mask = 16'h88A0;
defparam \Mux32~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N22
cycloneive_lcell_comb \Mux34~2 (
// Equation(s):
// \Mux34~2_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[26][29]~q ))) # (!temp_imemload_output_19 & (\storeregister[18][29]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[18][29]~q ),
	.datad(\storeregister[26][29]~q ),
	.cin(gnd),
	.combout(\Mux34~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~2 .lut_mask = 16'hDC98;
defparam \Mux34~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N2
cycloneive_lcell_comb \Mux34~4 (
// Equation(s):
// \Mux34~4_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18) # (\storeregister[24][29]~q )))) # (!temp_imemload_output_19 & (\storeregister[16][29]~q  & (!temp_imemload_output_18)))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[16][29]~q ),
	.datac(temp_imemload_output_18),
	.datad(\storeregister[24][29]~q ),
	.cin(gnd),
	.combout(\Mux34~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~4 .lut_mask = 16'hAEA4;
defparam \Mux34~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N2
cycloneive_lcell_comb \Mux34~12 (
// Equation(s):
// \Mux34~12_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][29]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & (\storeregister[4][29]~q )))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[4][29]~q ),
	.datad(\storeregister[5][29]~q ),
	.cin(gnd),
	.combout(\Mux34~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~12 .lut_mask = 16'hBA98;
defparam \Mux34~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N30
cycloneive_lcell_comb \Mux35~12 (
// Equation(s):
// \Mux35~12_combout  = (temp_imemload_output_17 & ((temp_imemload_output_16) # ((\storeregister[10][28]~q )))) # (!temp_imemload_output_17 & (!temp_imemload_output_16 & (\storeregister[8][28]~q )))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[8][28]~q ),
	.datad(\storeregister[10][28]~q ),
	.cin(gnd),
	.combout(\Mux35~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~12 .lut_mask = 16'hBA98;
defparam \Mux35~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N14
cycloneive_lcell_comb \Mux38~2 (
// Equation(s):
// \Mux38~2_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[26][25]~q ))) # (!temp_imemload_output_19 & (\storeregister[18][25]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[18][25]~q ),
	.datad(\storeregister[26][25]~q ),
	.cin(gnd),
	.combout(\Mux38~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~2 .lut_mask = 16'hDC98;
defparam \Mux38~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N30
cycloneive_lcell_comb \Mux38~12 (
// Equation(s):
// \Mux38~12_combout  = (temp_imemload_output_16 & ((\storeregister[5][25]~q ) # ((temp_imemload_output_17)))) # (!temp_imemload_output_16 & (((\storeregister[4][25]~q  & !temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[5][25]~q ),
	.datac(\storeregister[4][25]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux38~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~12 .lut_mask = 16'hAAD8;
defparam \Mux38~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N14
cycloneive_lcell_comb \Mux39~2 (
// Equation(s):
// \Mux39~2_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19) # (\storeregister[22][24]~q )))) # (!temp_imemload_output_18 & (\storeregister[18][24]~q  & (!temp_imemload_output_19)))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[18][24]~q ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[22][24]~q ),
	.cin(gnd),
	.combout(\Mux39~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~2 .lut_mask = 16'hAEA4;
defparam \Mux39~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N10
cycloneive_lcell_comb \Mux40~12 (
// Equation(s):
// \Mux40~12_combout  = (temp_imemload_output_16 & ((\storeregister[5][23]~q ) # ((temp_imemload_output_17)))) # (!temp_imemload_output_16 & (((\storeregister[4][23]~q  & !temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[5][23]~q ),
	.datac(\storeregister[4][23]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux40~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~12 .lut_mask = 16'hAAD8;
defparam \Mux40~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N26
cycloneive_lcell_comb \Mux42~2 (
// Equation(s):
// \Mux42~2_combout  = (temp_imemload_output_19 & ((\storeregister[26][21]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\storeregister[18][21]~q  & !temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[26][21]~q ),
	.datac(\storeregister[18][21]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux42~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~2 .lut_mask = 16'hAAD8;
defparam \Mux42~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N10
cycloneive_lcell_comb \Mux43~2 (
// Equation(s):
// \Mux43~2_combout  = (temp_imemload_output_18 & (((\storeregister[22][20]~q ) # (temp_imemload_output_19)))) # (!temp_imemload_output_18 & (\storeregister[18][20]~q  & ((!temp_imemload_output_19))))

	.dataa(\storeregister[18][20]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[22][20]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux43~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~2 .lut_mask = 16'hCCE2;
defparam \Mux43~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N16
cycloneive_lcell_comb \Mux49~4 (
// Equation(s):
// \Mux49~4_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[20][14]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[16][14]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[16][14]~q ),
	.datad(\storeregister[20][14]~q ),
	.cin(gnd),
	.combout(\Mux49~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~4 .lut_mask = 16'hBA98;
defparam \Mux49~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N14
cycloneive_lcell_comb \Mux54~2 (
// Equation(s):
// \Mux54~2_combout  = (temp_imemload_output_19 & ((\storeregister[26][9]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\storeregister[18][9]~q  & !temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[26][9]~q ),
	.datac(\storeregister[18][9]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux54~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~2 .lut_mask = 16'hAAD8;
defparam \Mux54~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N20
cycloneive_lcell_comb \Mux55~4 (
// Equation(s):
// \Mux55~4_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\storeregister[20][8]~q )) # (!temp_imemload_output_18 & ((\storeregister[16][8]~q )))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[20][8]~q ),
	.datac(\storeregister[16][8]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux55~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~4 .lut_mask = 16'hEE50;
defparam \Mux55~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N4
cycloneive_lcell_comb \Mux56~2 (
// Equation(s):
// \Mux56~2_combout  = (temp_imemload_output_19 & (((\storeregister[26][7]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[18][7]~q  & ((!temp_imemload_output_18))))

	.dataa(\storeregister[18][7]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[26][7]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux56~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~2 .lut_mask = 16'hCCE2;
defparam \Mux56~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N2
cycloneive_lcell_comb \Mux56~12 (
// Equation(s):
// \Mux56~12_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][7]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & (\storeregister[4][7]~q )))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[4][7]~q ),
	.datad(\storeregister[5][7]~q ),
	.cin(gnd),
	.combout(\Mux56~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~12 .lut_mask = 16'hBA98;
defparam \Mux56~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N18
cycloneive_lcell_comb \Mux57~4 (
// Equation(s):
// \Mux57~4_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[20][6]~q ))) # (!temp_imemload_output_18 & (\storeregister[16][6]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[16][6]~q ),
	.datac(temp_imemload_output_18),
	.datad(\storeregister[20][6]~q ),
	.cin(gnd),
	.combout(\Mux57~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~4 .lut_mask = 16'hF4A4;
defparam \Mux57~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N14
cycloneive_lcell_comb \Mux58~2 (
// Equation(s):
// \Mux58~2_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[26][5]~q ))) # (!temp_imemload_output_19 & (\storeregister[18][5]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[18][5]~q ),
	.datad(\storeregister[26][5]~q ),
	.cin(gnd),
	.combout(\Mux58~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~2 .lut_mask = 16'hDC98;
defparam \Mux58~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N12
cycloneive_lcell_comb \Mux50~2 (
// Equation(s):
// \Mux50~2_combout  = (temp_imemload_output_19 & (((\storeregister[26][13]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[18][13]~q  & ((!temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[18][13]~q ),
	.datac(\storeregister[26][13]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux50~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~2 .lut_mask = 16'hAAE4;
defparam \Mux50~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N30
cycloneive_lcell_comb \Mux52~14 (
// Equation(s):
// \Mux52~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][11]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][11]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[3][11]~q ),
	.datac(\storeregister[1][11]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux52~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~14 .lut_mask = 16'hD800;
defparam \Mux52~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N22
cycloneive_lcell_comb \Decoder0~13 (
// Equation(s):
// \Decoder0~13_combout  = (!temp_branchDest_01 & (temp_branchDest_11 & temp_regwrite2))

	.dataa(temp_branchDest_0),
	.datab(gnd),
	.datac(temp_branchDest_1),
	.datad(temp_regwrite),
	.cin(gnd),
	.combout(\Decoder0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~13 .lut_mask = 16'h5000;
defparam \Decoder0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N26
cycloneive_lcell_comb \Decoder0~20 (
// Equation(s):
// \Decoder0~20_combout  = (!temp_branchDest_01 & temp_regwrite2)

	.dataa(temp_branchDest_0),
	.datab(gnd),
	.datac(gnd),
	.datad(temp_regwrite),
	.cin(gnd),
	.combout(\Decoder0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~20 .lut_mask = 16'h5500;
defparam \Decoder0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N8
cycloneive_lcell_comb \storeregister[18][1]~feeder (
// Equation(s):
// \storeregister[18][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux30),
	.cin(gnd),
	.combout(\storeregister[18][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[18][1]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[18][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N6
cycloneive_lcell_comb \storeregister[28][2]~feeder (
// Equation(s):
// \storeregister[28][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux29),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[28][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][2]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[28][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N12
cycloneive_lcell_comb \storeregister[30][3]~feeder (
// Equation(s):
// \storeregister[30][3]~feeder_combout  = Mux28

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux28),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[30][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][3]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[30][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N12
cycloneive_lcell_comb \storeregister[20][13]~feeder (
// Equation(s):
// \storeregister[20][13]~feeder_combout  = Mux18

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux18),
	.cin(gnd),
	.combout(\storeregister[20][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][13]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[20][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N16
cycloneive_lcell_comb \storeregister[30][11]~feeder (
// Equation(s):
// \storeregister[30][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux20),
	.cin(gnd),
	.combout(\storeregister[30][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][11]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[30][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N2
cycloneive_lcell_comb \storeregister[18][31]~feeder (
// Equation(s):
// \storeregister[18][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux0),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[18][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[18][31]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[18][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N0
cycloneive_lcell_comb \storeregister[26][25]~feeder (
// Equation(s):
// \storeregister[26][25]~feeder_combout  = Mux6

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux6),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[26][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[26][25]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[26][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N12
cycloneive_lcell_comb \storeregister[28][28]~feeder (
// Equation(s):
// \storeregister[28][28]~feeder_combout  = Mux3

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux3),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[28][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][28]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[28][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N22
cycloneive_lcell_comb \storeregister[20][17]~feeder (
// Equation(s):
// \storeregister[20][17]~feeder_combout  = Mux14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux14),
	.cin(gnd),
	.combout(\storeregister[20][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][17]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[20][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N20
cycloneive_lcell_comb \storeregister[22][24]~feeder (
// Equation(s):
// \storeregister[22][24]~feeder_combout  = Mux7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux7),
	.cin(gnd),
	.combout(\storeregister[22][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[22][24]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[22][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N20
cycloneive_lcell_comb \storeregister[26][22]~feeder (
// Equation(s):
// \storeregister[26][22]~feeder_combout  = Mux9

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux9),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[26][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[26][22]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[26][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N26
cycloneive_lcell_comb \Mux62~9 (
// Equation(s):
// Mux62 = (temp_imemload_output_16 & ((\Mux62~6_combout  & (\Mux62~8_combout )) # (!\Mux62~6_combout  & ((\Mux62~1_combout ))))) # (!temp_imemload_output_16 & (((\Mux62~6_combout ))))

	.dataa(\Mux62~8_combout ),
	.datab(temp_imemload_output_16),
	.datac(\Mux62~1_combout ),
	.datad(\Mux62~6_combout ),
	.cin(gnd),
	.combout(Mux62),
	.cout());
// synopsys translate_off
defparam \Mux62~9 .lut_mask = 16'hBBC0;
defparam \Mux62~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N10
cycloneive_lcell_comb \Mux62~19 (
// Equation(s):
// Mux621 = (temp_imemload_output_18 & ((\Mux62~16_combout  & ((\Mux62~18_combout ))) # (!\Mux62~16_combout  & (\Mux62~11_combout )))) # (!temp_imemload_output_18 & (((\Mux62~16_combout ))))

	.dataa(\Mux62~11_combout ),
	.datab(temp_imemload_output_18),
	.datac(\Mux62~18_combout ),
	.datad(\Mux62~16_combout ),
	.cin(gnd),
	.combout(Mux621),
	.cout());
// synopsys translate_off
defparam \Mux62~19 .lut_mask = 16'hF388;
defparam \Mux62~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N6
cycloneive_lcell_comb \Mux30~9 (
// Equation(s):
// Mux301 = (temp_imemload_output_21 & ((\Mux30~6_combout  & ((\Mux30~8_combout ))) # (!\Mux30~6_combout  & (\Mux30~1_combout )))) # (!temp_imemload_output_21 & (\Mux30~6_combout ))

	.dataa(temp_imemload_output_21),
	.datab(\Mux30~6_combout ),
	.datac(\Mux30~1_combout ),
	.datad(\Mux30~8_combout ),
	.cin(gnd),
	.combout(Mux301),
	.cout());
// synopsys translate_off
defparam \Mux30~9 .lut_mask = 16'hEC64;
defparam \Mux30~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N2
cycloneive_lcell_comb \Mux30~19 (
// Equation(s):
// Mux302 = (\Mux30~16_combout  & (((\Mux30~18_combout ) # (!temp_imemload_output_23)))) # (!\Mux30~16_combout  & (\Mux30~11_combout  & (temp_imemload_output_23)))

	.dataa(\Mux30~11_combout ),
	.datab(\Mux30~16_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux30~18_combout ),
	.cin(gnd),
	.combout(Mux302),
	.cout());
// synopsys translate_off
defparam \Mux30~19 .lut_mask = 16'hEC2C;
defparam \Mux30~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N18
cycloneive_lcell_comb \Mux63~9 (
// Equation(s):
// Mux63 = (\Mux63~6_combout  & (((\Mux63~8_combout ) # (!temp_imemload_output_16)))) # (!\Mux63~6_combout  & (\Mux63~1_combout  & (temp_imemload_output_16)))

	.dataa(\Mux63~1_combout ),
	.datab(\Mux63~6_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux63~8_combout ),
	.cin(gnd),
	.combout(Mux63),
	.cout());
// synopsys translate_off
defparam \Mux63~9 .lut_mask = 16'hEC2C;
defparam \Mux63~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N10
cycloneive_lcell_comb \Mux63~19 (
// Equation(s):
// Mux631 = (temp_imemload_output_19 & ((\Mux63~16_combout  & ((\Mux63~18_combout ))) # (!\Mux63~16_combout  & (\Mux63~11_combout )))) # (!temp_imemload_output_19 & (((\Mux63~16_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\Mux63~11_combout ),
	.datac(\Mux63~16_combout ),
	.datad(\Mux63~18_combout ),
	.cin(gnd),
	.combout(Mux631),
	.cout());
// synopsys translate_off
defparam \Mux63~19 .lut_mask = 16'hF858;
defparam \Mux63~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N16
cycloneive_lcell_comb \Mux31~9 (
// Equation(s):
// Mux311 = (temp_imemload_output_21 & ((\Mux31~6_combout  & ((\Mux31~8_combout ))) # (!\Mux31~6_combout  & (\Mux31~1_combout )))) # (!temp_imemload_output_21 & (((\Mux31~6_combout ))))

	.dataa(\Mux31~1_combout ),
	.datab(\Mux31~8_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux31~6_combout ),
	.cin(gnd),
	.combout(Mux311),
	.cout());
// synopsys translate_off
defparam \Mux31~9 .lut_mask = 16'hCFA0;
defparam \Mux31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N26
cycloneive_lcell_comb \Mux31~19 (
// Equation(s):
// Mux312 = (\Mux31~16_combout  & (((\Mux31~18_combout ) # (!temp_imemload_output_24)))) # (!\Mux31~16_combout  & (\Mux31~11_combout  & ((temp_imemload_output_24))))

	.dataa(\Mux31~16_combout ),
	.datab(\Mux31~11_combout ),
	.datac(\Mux31~18_combout ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(Mux312),
	.cout());
// synopsys translate_off
defparam \Mux31~19 .lut_mask = 16'hE4AA;
defparam \Mux31~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N20
cycloneive_lcell_comb \Mux29~9 (
// Equation(s):
// Mux291 = (\Mux29~6_combout  & (((\Mux29~8_combout )) # (!temp_imemload_output_21))) # (!\Mux29~6_combout  & (temp_imemload_output_21 & ((\Mux29~1_combout ))))

	.dataa(\Mux29~6_combout ),
	.datab(temp_imemload_output_21),
	.datac(\Mux29~8_combout ),
	.datad(\Mux29~1_combout ),
	.cin(gnd),
	.combout(Mux291),
	.cout());
// synopsys translate_off
defparam \Mux29~9 .lut_mask = 16'hE6A2;
defparam \Mux29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N14
cycloneive_lcell_comb \Mux29~19 (
// Equation(s):
// Mux292 = (\Mux29~16_combout  & (((\Mux29~18_combout )) # (!temp_imemload_output_24))) # (!\Mux29~16_combout  & (temp_imemload_output_24 & ((\Mux29~11_combout ))))

	.dataa(\Mux29~16_combout ),
	.datab(temp_imemload_output_24),
	.datac(\Mux29~18_combout ),
	.datad(\Mux29~11_combout ),
	.cin(gnd),
	.combout(Mux292),
	.cout());
// synopsys translate_off
defparam \Mux29~19 .lut_mask = 16'hE6A2;
defparam \Mux29~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N10
cycloneive_lcell_comb \Mux27~9 (
// Equation(s):
// Mux271 = (\Mux27~6_combout  & ((\Mux27~8_combout ) # ((!temp_imemload_output_21)))) # (!\Mux27~6_combout  & (((temp_imemload_output_21 & \Mux27~1_combout ))))

	.dataa(\Mux27~8_combout ),
	.datab(\Mux27~6_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux27~1_combout ),
	.cin(gnd),
	.combout(Mux271),
	.cout());
// synopsys translate_off
defparam \Mux27~9 .lut_mask = 16'hBC8C;
defparam \Mux27~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N16
cycloneive_lcell_comb \Mux27~19 (
// Equation(s):
// Mux272 = (\Mux27~16_combout  & (((\Mux27~18_combout ) # (!temp_imemload_output_24)))) # (!\Mux27~16_combout  & (\Mux27~11_combout  & (temp_imemload_output_24)))

	.dataa(\Mux27~16_combout ),
	.datab(\Mux27~11_combout ),
	.datac(temp_imemload_output_24),
	.datad(\Mux27~18_combout ),
	.cin(gnd),
	.combout(Mux272),
	.cout());
// synopsys translate_off
defparam \Mux27~19 .lut_mask = 16'hEA4A;
defparam \Mux27~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N20
cycloneive_lcell_comb \Mux28~9 (
// Equation(s):
// Mux281 = (\Mux28~6_combout  & (((\Mux28~8_combout ) # (!temp_imemload_output_21)))) # (!\Mux28~6_combout  & (\Mux28~1_combout  & (temp_imemload_output_21)))

	.dataa(\Mux28~6_combout ),
	.datab(\Mux28~1_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux28~8_combout ),
	.cin(gnd),
	.combout(Mux281),
	.cout());
// synopsys translate_off
defparam \Mux28~9 .lut_mask = 16'hEA4A;
defparam \Mux28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N18
cycloneive_lcell_comb \Mux28~19 (
// Equation(s):
// Mux282 = (\Mux28~16_combout  & (((\Mux28~18_combout ) # (!temp_imemload_output_23)))) # (!\Mux28~16_combout  & (\Mux28~11_combout  & (temp_imemload_output_23)))

	.dataa(\Mux28~11_combout ),
	.datab(\Mux28~16_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux28~18_combout ),
	.cin(gnd),
	.combout(Mux282),
	.cout());
// synopsys translate_off
defparam \Mux28~19 .lut_mask = 16'hEC2C;
defparam \Mux28~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N14
cycloneive_lcell_comb \Mux61~9 (
// Equation(s):
// Mux61 = (\Mux61~6_combout  & (((\Mux61~8_combout ) # (!temp_imemload_output_16)))) # (!\Mux61~6_combout  & (\Mux61~1_combout  & (temp_imemload_output_16)))

	.dataa(\Mux61~6_combout ),
	.datab(\Mux61~1_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux61~8_combout ),
	.cin(gnd),
	.combout(Mux61),
	.cout());
// synopsys translate_off
defparam \Mux61~9 .lut_mask = 16'hEA4A;
defparam \Mux61~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N12
cycloneive_lcell_comb \Mux61~19 (
// Equation(s):
// Mux611 = (temp_imemload_output_18 & ((\Mux61~16_combout  & ((\Mux61~18_combout ))) # (!\Mux61~16_combout  & (\Mux61~11_combout )))) # (!temp_imemload_output_18 & (\Mux61~16_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux61~16_combout ),
	.datac(\Mux61~11_combout ),
	.datad(\Mux61~18_combout ),
	.cin(gnd),
	.combout(Mux611),
	.cout());
// synopsys translate_off
defparam \Mux61~19 .lut_mask = 16'hEC64;
defparam \Mux61~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N16
cycloneive_lcell_comb \Mux23~9 (
// Equation(s):
// Mux231 = (temp_imemload_output_21 & ((\Mux23~6_combout  & (\Mux23~8_combout )) # (!\Mux23~6_combout  & ((\Mux23~1_combout ))))) # (!temp_imemload_output_21 & (((\Mux23~6_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux23~8_combout ),
	.datac(\Mux23~6_combout ),
	.datad(\Mux23~1_combout ),
	.cin(gnd),
	.combout(Mux231),
	.cout());
// synopsys translate_off
defparam \Mux23~9 .lut_mask = 16'hDAD0;
defparam \Mux23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N4
cycloneive_lcell_comb \Mux23~19 (
// Equation(s):
// Mux232 = (temp_imemload_output_24 & ((\Mux23~16_combout  & ((\Mux23~18_combout ))) # (!\Mux23~16_combout  & (\Mux23~11_combout )))) # (!temp_imemload_output_24 & (((\Mux23~16_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\Mux23~11_combout ),
	.datac(\Mux23~16_combout ),
	.datad(\Mux23~18_combout ),
	.cin(gnd),
	.combout(Mux232),
	.cout());
// synopsys translate_off
defparam \Mux23~19 .lut_mask = 16'hF858;
defparam \Mux23~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N26
cycloneive_lcell_comb \Mux24~9 (
// Equation(s):
// Mux241 = (temp_imemload_output_21 & ((\Mux24~6_combout  & ((\Mux24~8_combout ))) # (!\Mux24~6_combout  & (\Mux24~1_combout )))) # (!temp_imemload_output_21 & (((\Mux24~6_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux24~1_combout ),
	.datac(\Mux24~8_combout ),
	.datad(\Mux24~6_combout ),
	.cin(gnd),
	.combout(Mux241),
	.cout());
// synopsys translate_off
defparam \Mux24~9 .lut_mask = 16'hF588;
defparam \Mux24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N30
cycloneive_lcell_comb \Mux24~19 (
// Equation(s):
// Mux242 = (temp_imemload_output_23 & ((\Mux24~16_combout  & ((\Mux24~18_combout ))) # (!\Mux24~16_combout  & (\Mux24~11_combout )))) # (!temp_imemload_output_23 & (((\Mux24~16_combout ))))

	.dataa(\Mux24~11_combout ),
	.datab(temp_imemload_output_23),
	.datac(\Mux24~18_combout ),
	.datad(\Mux24~16_combout ),
	.cin(gnd),
	.combout(Mux242),
	.cout());
// synopsys translate_off
defparam \Mux24~19 .lut_mask = 16'hF388;
defparam \Mux24~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N16
cycloneive_lcell_comb \Mux25~9 (
// Equation(s):
// Mux251 = (\Mux25~6_combout  & ((\Mux25~8_combout ) # ((!temp_imemload_output_21)))) # (!\Mux25~6_combout  & (((\Mux25~1_combout  & temp_imemload_output_21))))

	.dataa(\Mux25~6_combout ),
	.datab(\Mux25~8_combout ),
	.datac(\Mux25~1_combout ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(Mux251),
	.cout());
// synopsys translate_off
defparam \Mux25~9 .lut_mask = 16'hD8AA;
defparam \Mux25~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N16
cycloneive_lcell_comb \Mux25~19 (
// Equation(s):
// Mux252 = (temp_imemload_output_24 & ((\Mux25~16_combout  & ((\Mux25~18_combout ))) # (!\Mux25~16_combout  & (\Mux25~11_combout )))) # (!temp_imemload_output_24 & (((\Mux25~16_combout ))))

	.dataa(\Mux25~11_combout ),
	.datab(temp_imemload_output_24),
	.datac(\Mux25~16_combout ),
	.datad(\Mux25~18_combout ),
	.cin(gnd),
	.combout(Mux252),
	.cout());
// synopsys translate_off
defparam \Mux25~19 .lut_mask = 16'hF838;
defparam \Mux25~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N12
cycloneive_lcell_comb \Mux26~9 (
// Equation(s):
// Mux261 = (\Mux26~6_combout  & ((\Mux26~8_combout ) # ((!temp_imemload_output_21)))) # (!\Mux26~6_combout  & (((temp_imemload_output_21 & \Mux26~1_combout ))))

	.dataa(\Mux26~6_combout ),
	.datab(\Mux26~8_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux26~1_combout ),
	.cin(gnd),
	.combout(Mux261),
	.cout());
// synopsys translate_off
defparam \Mux26~9 .lut_mask = 16'hDA8A;
defparam \Mux26~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N24
cycloneive_lcell_comb \Mux26~19 (
// Equation(s):
// Mux262 = (temp_imemload_output_23 & ((\Mux26~16_combout  & (\Mux26~18_combout )) # (!\Mux26~16_combout  & ((\Mux26~11_combout ))))) # (!temp_imemload_output_23 & (\Mux26~16_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux26~16_combout ),
	.datac(\Mux26~18_combout ),
	.datad(\Mux26~11_combout ),
	.cin(gnd),
	.combout(Mux262),
	.cout());
// synopsys translate_off
defparam \Mux26~19 .lut_mask = 16'hE6C4;
defparam \Mux26~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N2
cycloneive_lcell_comb \Mux60~9 (
// Equation(s):
// Mux60 = (temp_imemload_output_16 & ((\Mux60~6_combout  & ((\Mux60~8_combout ))) # (!\Mux60~6_combout  & (\Mux60~1_combout )))) # (!temp_imemload_output_16 & (\Mux60~6_combout ))

	.dataa(temp_imemload_output_16),
	.datab(\Mux60~6_combout ),
	.datac(\Mux60~1_combout ),
	.datad(\Mux60~8_combout ),
	.cin(gnd),
	.combout(Mux60),
	.cout());
// synopsys translate_off
defparam \Mux60~9 .lut_mask = 16'hEC64;
defparam \Mux60~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N2
cycloneive_lcell_comb \Mux60~19 (
// Equation(s):
// Mux601 = (\Mux60~16_combout  & ((\Mux60~18_combout ) # ((!temp_imemload_output_19)))) # (!\Mux60~16_combout  & (((\Mux60~11_combout  & temp_imemload_output_19))))

	.dataa(\Mux60~16_combout ),
	.datab(\Mux60~18_combout ),
	.datac(\Mux60~11_combout ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(Mux601),
	.cout());
// synopsys translate_off
defparam \Mux60~19 .lut_mask = 16'hD8AA;
defparam \Mux60~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N14
cycloneive_lcell_comb \Mux15~9 (
// Equation(s):
// Mux151 = (\Mux15~6_combout  & (((\Mux15~8_combout ) # (!temp_imemload_output_21)))) # (!\Mux15~6_combout  & (\Mux15~1_combout  & ((temp_imemload_output_21))))

	.dataa(\Mux15~1_combout ),
	.datab(\Mux15~6_combout ),
	.datac(\Mux15~8_combout ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(Mux151),
	.cout());
// synopsys translate_off
defparam \Mux15~9 .lut_mask = 16'hE2CC;
defparam \Mux15~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N4
cycloneive_lcell_comb \Mux15~19 (
// Equation(s):
// Mux152 = (temp_imemload_output_24 & ((\Mux15~16_combout  & ((\Mux15~18_combout ))) # (!\Mux15~16_combout  & (\Mux15~11_combout )))) # (!temp_imemload_output_24 & (((\Mux15~16_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\Mux15~11_combout ),
	.datac(\Mux15~16_combout ),
	.datad(\Mux15~18_combout ),
	.cin(gnd),
	.combout(Mux152),
	.cout());
// synopsys translate_off
defparam \Mux15~19 .lut_mask = 16'hF858;
defparam \Mux15~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N14
cycloneive_lcell_comb \Mux17~9 (
// Equation(s):
// Mux171 = (\Mux17~6_combout  & ((\Mux17~8_combout ) # ((!temp_imemload_output_21)))) # (!\Mux17~6_combout  & (((temp_imemload_output_21 & \Mux17~1_combout ))))

	.dataa(\Mux17~8_combout ),
	.datab(\Mux17~6_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux17~1_combout ),
	.cin(gnd),
	.combout(Mux171),
	.cout());
// synopsys translate_off
defparam \Mux17~9 .lut_mask = 16'hBC8C;
defparam \Mux17~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N12
cycloneive_lcell_comb \Mux17~19 (
// Equation(s):
// Mux172 = (temp_imemload_output_24 & ((\Mux17~16_combout  & (\Mux17~18_combout )) # (!\Mux17~16_combout  & ((\Mux17~11_combout ))))) # (!temp_imemload_output_24 & (((\Mux17~16_combout ))))

	.dataa(\Mux17~18_combout ),
	.datab(temp_imemload_output_24),
	.datac(\Mux17~11_combout ),
	.datad(\Mux17~16_combout ),
	.cin(gnd),
	.combout(Mux172),
	.cout());
// synopsys translate_off
defparam \Mux17~19 .lut_mask = 16'hBBC0;
defparam \Mux17~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N20
cycloneive_lcell_comb \Mux16~9 (
// Equation(s):
// Mux161 = (\Mux16~6_combout  & (((\Mux16~8_combout ) # (!temp_imemload_output_21)))) # (!\Mux16~6_combout  & (\Mux16~1_combout  & (temp_imemload_output_21)))

	.dataa(\Mux16~6_combout ),
	.datab(\Mux16~1_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux16~8_combout ),
	.cin(gnd),
	.combout(Mux161),
	.cout());
// synopsys translate_off
defparam \Mux16~9 .lut_mask = 16'hEA4A;
defparam \Mux16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N28
cycloneive_lcell_comb \Mux16~19 (
// Equation(s):
// Mux162 = (temp_imemload_output_23 & ((\Mux16~16_combout  & ((\Mux16~18_combout ))) # (!\Mux16~16_combout  & (\Mux16~11_combout )))) # (!temp_imemload_output_23 & (((\Mux16~16_combout ))))

	.dataa(\Mux16~11_combout ),
	.datab(temp_imemload_output_23),
	.datac(\Mux16~18_combout ),
	.datad(\Mux16~16_combout ),
	.cin(gnd),
	.combout(Mux162),
	.cout());
// synopsys translate_off
defparam \Mux16~19 .lut_mask = 16'hF388;
defparam \Mux16~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N14
cycloneive_lcell_comb \Mux18~9 (
// Equation(s):
// Mux181 = (\Mux18~6_combout  & ((\Mux18~8_combout ) # ((!temp_imemload_output_21)))) # (!\Mux18~6_combout  & (((\Mux18~1_combout  & temp_imemload_output_21))))

	.dataa(\Mux18~8_combout ),
	.datab(\Mux18~1_combout ),
	.datac(\Mux18~6_combout ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(Mux181),
	.cout());
// synopsys translate_off
defparam \Mux18~9 .lut_mask = 16'hACF0;
defparam \Mux18~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N16
cycloneive_lcell_comb \Mux18~19 (
// Equation(s):
// Mux182 = (\Mux18~16_combout  & (((\Mux18~18_combout ) # (!temp_imemload_output_23)))) # (!\Mux18~16_combout  & (\Mux18~11_combout  & (temp_imemload_output_23)))

	.dataa(\Mux18~16_combout ),
	.datab(\Mux18~11_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux18~18_combout ),
	.cin(gnd),
	.combout(Mux182),
	.cout());
// synopsys translate_off
defparam \Mux18~19 .lut_mask = 16'hEA4A;
defparam \Mux18~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N6
cycloneive_lcell_comb \Mux19~9 (
// Equation(s):
// Mux191 = (temp_imemload_output_21 & ((\Mux19~6_combout  & ((\Mux19~8_combout ))) # (!\Mux19~6_combout  & (\Mux19~1_combout )))) # (!temp_imemload_output_21 & (((\Mux19~6_combout ))))

	.dataa(\Mux19~1_combout ),
	.datab(temp_imemload_output_21),
	.datac(\Mux19~6_combout ),
	.datad(\Mux19~8_combout ),
	.cin(gnd),
	.combout(Mux191),
	.cout());
// synopsys translate_off
defparam \Mux19~9 .lut_mask = 16'hF838;
defparam \Mux19~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N18
cycloneive_lcell_comb \Mux19~19 (
// Equation(s):
// Mux192 = (\Mux19~16_combout  & (((\Mux19~18_combout )) # (!temp_imemload_output_24))) # (!\Mux19~16_combout  & (temp_imemload_output_24 & ((\Mux19~11_combout ))))

	.dataa(\Mux19~16_combout ),
	.datab(temp_imemload_output_24),
	.datac(\Mux19~18_combout ),
	.datad(\Mux19~11_combout ),
	.cin(gnd),
	.combout(Mux192),
	.cout());
// synopsys translate_off
defparam \Mux19~19 .lut_mask = 16'hE6A2;
defparam \Mux19~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N18
cycloneive_lcell_comb \Mux21~9 (
// Equation(s):
// Mux211 = (temp_imemload_output_21 & ((\Mux21~6_combout  & ((\Mux21~8_combout ))) # (!\Mux21~6_combout  & (\Mux21~1_combout )))) # (!temp_imemload_output_21 & (\Mux21~6_combout ))

	.dataa(temp_imemload_output_21),
	.datab(\Mux21~6_combout ),
	.datac(\Mux21~1_combout ),
	.datad(\Mux21~8_combout ),
	.cin(gnd),
	.combout(Mux211),
	.cout());
// synopsys translate_off
defparam \Mux21~9 .lut_mask = 16'hEC64;
defparam \Mux21~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N18
cycloneive_lcell_comb \Mux21~19 (
// Equation(s):
// Mux212 = (temp_imemload_output_24 & ((\Mux21~16_combout  & ((\Mux21~18_combout ))) # (!\Mux21~16_combout  & (\Mux21~11_combout )))) # (!temp_imemload_output_24 & (((\Mux21~16_combout ))))

	.dataa(\Mux21~11_combout ),
	.datab(temp_imemload_output_24),
	.datac(\Mux21~16_combout ),
	.datad(\Mux21~18_combout ),
	.cin(gnd),
	.combout(Mux212),
	.cout());
// synopsys translate_off
defparam \Mux21~19 .lut_mask = 16'hF838;
defparam \Mux21~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N16
cycloneive_lcell_comb \Mux20~9 (
// Equation(s):
// Mux201 = (\Mux20~6_combout  & (((\Mux20~8_combout ) # (!temp_imemload_output_21)))) # (!\Mux20~6_combout  & (\Mux20~1_combout  & (temp_imemload_output_21)))

	.dataa(\Mux20~6_combout ),
	.datab(\Mux20~1_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux20~8_combout ),
	.cin(gnd),
	.combout(Mux201),
	.cout());
// synopsys translate_off
defparam \Mux20~9 .lut_mask = 16'hEA4A;
defparam \Mux20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N20
cycloneive_lcell_comb \Mux20~19 (
// Equation(s):
// Mux202 = (\Mux20~16_combout  & (((\Mux20~18_combout ) # (!temp_imemload_output_23)))) # (!\Mux20~16_combout  & (\Mux20~11_combout  & (temp_imemload_output_23)))

	.dataa(\Mux20~11_combout ),
	.datab(\Mux20~16_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux20~18_combout ),
	.cin(gnd),
	.combout(Mux202),
	.cout());
// synopsys translate_off
defparam \Mux20~19 .lut_mask = 16'hEC2C;
defparam \Mux20~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N0
cycloneive_lcell_comb \Mux22~9 (
// Equation(s):
// Mux221 = (temp_imemload_output_21 & ((\Mux22~6_combout  & ((\Mux22~8_combout ))) # (!\Mux22~6_combout  & (\Mux22~1_combout )))) # (!temp_imemload_output_21 & (((\Mux22~6_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux22~1_combout ),
	.datac(\Mux22~6_combout ),
	.datad(\Mux22~8_combout ),
	.cin(gnd),
	.combout(Mux221),
	.cout());
// synopsys translate_off
defparam \Mux22~9 .lut_mask = 16'hF858;
defparam \Mux22~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N16
cycloneive_lcell_comb \Mux22~19 (
// Equation(s):
// Mux222 = (temp_imemload_output_23 & ((\Mux22~16_combout  & ((\Mux22~18_combout ))) # (!\Mux22~16_combout  & (\Mux22~11_combout )))) # (!temp_imemload_output_23 & (((\Mux22~16_combout ))))

	.dataa(\Mux22~11_combout ),
	.datab(\Mux22~18_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux22~16_combout ),
	.cin(gnd),
	.combout(Mux222),
	.cout());
// synopsys translate_off
defparam \Mux22~19 .lut_mask = 16'hCFA0;
defparam \Mux22~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N16
cycloneive_lcell_comb \Mux59~9 (
// Equation(s):
// Mux59 = (\Mux59~6_combout  & ((\Mux59~8_combout ) # ((!temp_imemload_output_16)))) # (!\Mux59~6_combout  & (((\Mux59~1_combout  & temp_imemload_output_16))))

	.dataa(\Mux59~8_combout ),
	.datab(\Mux59~1_combout ),
	.datac(\Mux59~6_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(Mux59),
	.cout());
// synopsys translate_off
defparam \Mux59~9 .lut_mask = 16'hACF0;
defparam \Mux59~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N28
cycloneive_lcell_comb \Mux59~19 (
// Equation(s):
// Mux591 = (\Mux59~16_combout  & ((\Mux59~18_combout ) # ((!temp_imemload_output_18)))) # (!\Mux59~16_combout  & (((\Mux59~11_combout  & temp_imemload_output_18))))

	.dataa(\Mux59~16_combout ),
	.datab(\Mux59~18_combout ),
	.datac(\Mux59~11_combout ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(Mux591),
	.cout());
// synopsys translate_off
defparam \Mux59~19 .lut_mask = 16'hD8AA;
defparam \Mux59~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N26
cycloneive_lcell_comb \Mux0~9 (
// Equation(s):
// Mux01 = (\Mux0~6_combout  & ((\Mux0~8_combout ) # ((!temp_imemload_output_21)))) # (!\Mux0~6_combout  & (((\Mux0~1_combout  & temp_imemload_output_21))))

	.dataa(\Mux0~8_combout ),
	.datab(\Mux0~6_combout ),
	.datac(\Mux0~1_combout ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(Mux01),
	.cout());
// synopsys translate_off
defparam \Mux0~9 .lut_mask = 16'hB8CC;
defparam \Mux0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N10
cycloneive_lcell_comb \Mux0~19 (
// Equation(s):
// Mux02 = (\Mux0~16_combout  & ((\Mux0~18_combout ) # ((!temp_imemload_output_23)))) # (!\Mux0~16_combout  & (((\Mux0~11_combout  & temp_imemload_output_23))))

	.dataa(\Mux0~18_combout ),
	.datab(\Mux0~16_combout ),
	.datac(\Mux0~11_combout ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(Mux02),
	.cout());
// synopsys translate_off
defparam \Mux0~19 .lut_mask = 16'hB8CC;
defparam \Mux0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N22
cycloneive_lcell_comb \Mux1~9 (
// Equation(s):
// Mux110 = (\Mux1~6_combout  & (((\Mux1~8_combout ) # (!temp_imemload_output_21)))) # (!\Mux1~6_combout  & (\Mux1~1_combout  & (temp_imemload_output_21)))

	.dataa(\Mux1~1_combout ),
	.datab(\Mux1~6_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux1~8_combout ),
	.cin(gnd),
	.combout(Mux110),
	.cout());
// synopsys translate_off
defparam \Mux1~9 .lut_mask = 16'hEC2C;
defparam \Mux1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N6
cycloneive_lcell_comb \Mux1~19 (
// Equation(s):
// Mux111 = (temp_imemload_output_24 & ((\Mux1~16_combout  & (\Mux1~18_combout )) # (!\Mux1~16_combout  & ((\Mux1~11_combout ))))) # (!temp_imemload_output_24 & (((\Mux1~16_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\Mux1~18_combout ),
	.datac(\Mux1~16_combout ),
	.datad(\Mux1~11_combout ),
	.cin(gnd),
	.combout(Mux111),
	.cout());
// synopsys translate_off
defparam \Mux1~19 .lut_mask = 16'hDAD0;
defparam \Mux1~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N14
cycloneive_lcell_comb \Mux2~9 (
// Equation(s):
// Mux210 = (\Mux2~6_combout  & (((\Mux2~8_combout ) # (!temp_imemload_output_21)))) # (!\Mux2~6_combout  & (\Mux2~1_combout  & (temp_imemload_output_21)))

	.dataa(\Mux2~6_combout ),
	.datab(\Mux2~1_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux2~8_combout ),
	.cin(gnd),
	.combout(Mux210),
	.cout());
// synopsys translate_off
defparam \Mux2~9 .lut_mask = 16'hEA4A;
defparam \Mux2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N20
cycloneive_lcell_comb \Mux2~19 (
// Equation(s):
// Mux213 = (\Mux2~16_combout  & ((\Mux2~18_combout ) # ((!temp_imemload_output_23)))) # (!\Mux2~16_combout  & (((temp_imemload_output_23 & \Mux2~11_combout ))))

	.dataa(\Mux2~18_combout ),
	.datab(\Mux2~16_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux2~11_combout ),
	.cin(gnd),
	.combout(Mux213),
	.cout());
// synopsys translate_off
defparam \Mux2~19 .lut_mask = 16'hBC8C;
defparam \Mux2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N4
cycloneive_lcell_comb \Mux5~9 (
// Equation(s):
// Mux51 = (temp_imemload_output_21 & ((\Mux5~6_combout  & (\Mux5~8_combout )) # (!\Mux5~6_combout  & ((\Mux5~1_combout ))))) # (!temp_imemload_output_21 & (((\Mux5~6_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux5~8_combout ),
	.datac(\Mux5~6_combout ),
	.datad(\Mux5~1_combout ),
	.cin(gnd),
	.combout(Mux51),
	.cout());
// synopsys translate_off
defparam \Mux5~9 .lut_mask = 16'hDAD0;
defparam \Mux5~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N18
cycloneive_lcell_comb \Mux5~19 (
// Equation(s):
// Mux52 = (temp_imemload_output_24 & ((\Mux5~16_combout  & ((\Mux5~18_combout ))) # (!\Mux5~16_combout  & (\Mux5~11_combout )))) # (!temp_imemload_output_24 & (((\Mux5~16_combout ))))

	.dataa(\Mux5~11_combout ),
	.datab(\Mux5~18_combout ),
	.datac(temp_imemload_output_24),
	.datad(\Mux5~16_combout ),
	.cin(gnd),
	.combout(Mux52),
	.cout());
// synopsys translate_off
defparam \Mux5~19 .lut_mask = 16'hCFA0;
defparam \Mux5~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N22
cycloneive_lcell_comb \Mux6~9 (
// Equation(s):
// Mux64 = (\Mux6~6_combout  & ((\Mux6~8_combout ) # ((!temp_imemload_output_21)))) # (!\Mux6~6_combout  & (((temp_imemload_output_21 & \Mux6~1_combout ))))

	.dataa(\Mux6~6_combout ),
	.datab(\Mux6~8_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux6~1_combout ),
	.cin(gnd),
	.combout(Mux64),
	.cout());
// synopsys translate_off
defparam \Mux6~9 .lut_mask = 16'hDA8A;
defparam \Mux6~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N22
cycloneive_lcell_comb \Mux6~19 (
// Equation(s):
// Mux65 = (temp_imemload_output_23 & ((\Mux6~16_combout  & (\Mux6~18_combout )) # (!\Mux6~16_combout  & ((\Mux6~11_combout ))))) # (!temp_imemload_output_23 & (((\Mux6~16_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\Mux6~18_combout ),
	.datac(\Mux6~16_combout ),
	.datad(\Mux6~11_combout ),
	.cin(gnd),
	.combout(Mux65),
	.cout());
// synopsys translate_off
defparam \Mux6~19 .lut_mask = 16'hDAD0;
defparam \Mux6~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N24
cycloneive_lcell_comb \Mux3~9 (
// Equation(s):
// Mux32 = (temp_imemload_output_21 & ((\Mux3~6_combout  & (\Mux3~8_combout )) # (!\Mux3~6_combout  & ((\Mux3~1_combout ))))) # (!temp_imemload_output_21 & (\Mux3~6_combout ))

	.dataa(temp_imemload_output_21),
	.datab(\Mux3~6_combout ),
	.datac(\Mux3~8_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(Mux32),
	.cout());
// synopsys translate_off
defparam \Mux3~9 .lut_mask = 16'hE6C4;
defparam \Mux3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y40_N30
cycloneive_lcell_comb \Mux3~19 (
// Equation(s):
// Mux33 = (temp_imemload_output_24 & ((\Mux3~16_combout  & ((\Mux3~18_combout ))) # (!\Mux3~16_combout  & (\Mux3~11_combout )))) # (!temp_imemload_output_24 & (((\Mux3~16_combout ))))

	.dataa(\Mux3~11_combout ),
	.datab(\Mux3~18_combout ),
	.datac(temp_imemload_output_24),
	.datad(\Mux3~16_combout ),
	.cin(gnd),
	.combout(Mux33),
	.cout());
// synopsys translate_off
defparam \Mux3~19 .lut_mask = 16'hCFA0;
defparam \Mux3~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N10
cycloneive_lcell_comb \Mux4~9 (
// Equation(s):
// Mux41 = (temp_imemload_output_21 & ((\Mux4~6_combout  & (\Mux4~8_combout )) # (!\Mux4~6_combout  & ((\Mux4~1_combout ))))) # (!temp_imemload_output_21 & (((\Mux4~6_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux4~8_combout ),
	.datac(\Mux4~1_combout ),
	.datad(\Mux4~6_combout ),
	.cin(gnd),
	.combout(Mux41),
	.cout());
// synopsys translate_off
defparam \Mux4~9 .lut_mask = 16'hDDA0;
defparam \Mux4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N14
cycloneive_lcell_comb \Mux4~19 (
// Equation(s):
// Mux42 = (temp_imemload_output_23 & ((\Mux4~16_combout  & ((\Mux4~18_combout ))) # (!\Mux4~16_combout  & (\Mux4~11_combout )))) # (!temp_imemload_output_23 & (((\Mux4~16_combout ))))

	.dataa(\Mux4~11_combout ),
	.datab(temp_imemload_output_23),
	.datac(\Mux4~16_combout ),
	.datad(\Mux4~18_combout ),
	.cin(gnd),
	.combout(Mux42),
	.cout());
// synopsys translate_off
defparam \Mux4~19 .lut_mask = 16'hF838;
defparam \Mux4~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N6
cycloneive_lcell_comb \Mux14~9 (
// Equation(s):
// Mux141 = (\Mux14~6_combout  & ((\Mux14~8_combout ) # ((!temp_imemload_output_21)))) # (!\Mux14~6_combout  & (((temp_imemload_output_21 & \Mux14~1_combout ))))

	.dataa(\Mux14~6_combout ),
	.datab(\Mux14~8_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux14~1_combout ),
	.cin(gnd),
	.combout(Mux141),
	.cout());
// synopsys translate_off
defparam \Mux14~9 .lut_mask = 16'hDA8A;
defparam \Mux14~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N20
cycloneive_lcell_comb \Mux14~19 (
// Equation(s):
// Mux142 = (\Mux14~16_combout  & ((\Mux14~18_combout ) # ((!temp_imemload_output_23)))) # (!\Mux14~16_combout  & (((temp_imemload_output_23 & \Mux14~11_combout ))))

	.dataa(\Mux14~18_combout ),
	.datab(\Mux14~16_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux14~11_combout ),
	.cin(gnd),
	.combout(Mux142),
	.cout());
// synopsys translate_off
defparam \Mux14~19 .lut_mask = 16'hBC8C;
defparam \Mux14~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N22
cycloneive_lcell_comb \Mux11~9 (
// Equation(s):
// Mux112 = (temp_imemload_output_21 & ((\Mux11~6_combout  & (\Mux11~8_combout )) # (!\Mux11~6_combout  & ((\Mux11~1_combout ))))) # (!temp_imemload_output_21 & (((\Mux11~6_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux11~8_combout ),
	.datac(\Mux11~1_combout ),
	.datad(\Mux11~6_combout ),
	.cin(gnd),
	.combout(Mux112),
	.cout());
// synopsys translate_off
defparam \Mux11~9 .lut_mask = 16'hDDA0;
defparam \Mux11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N18
cycloneive_lcell_comb \Mux11~19 (
// Equation(s):
// Mux113 = (temp_imemload_output_24 & ((\Mux11~16_combout  & (\Mux11~18_combout )) # (!\Mux11~16_combout  & ((\Mux11~11_combout ))))) # (!temp_imemload_output_24 & (((\Mux11~16_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\Mux11~18_combout ),
	.datac(\Mux11~16_combout ),
	.datad(\Mux11~11_combout ),
	.cin(gnd),
	.combout(Mux113),
	.cout());
// synopsys translate_off
defparam \Mux11~19 .lut_mask = 16'hDAD0;
defparam \Mux11~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N8
cycloneive_lcell_comb \Mux12~9 (
// Equation(s):
// Mux121 = (temp_imemload_output_21 & ((\Mux12~6_combout  & ((\Mux12~8_combout ))) # (!\Mux12~6_combout  & (\Mux12~1_combout )))) # (!temp_imemload_output_21 & (\Mux12~6_combout ))

	.dataa(temp_imemload_output_21),
	.datab(\Mux12~6_combout ),
	.datac(\Mux12~1_combout ),
	.datad(\Mux12~8_combout ),
	.cin(gnd),
	.combout(Mux121),
	.cout());
// synopsys translate_off
defparam \Mux12~9 .lut_mask = 16'hEC64;
defparam \Mux12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N28
cycloneive_lcell_comb \Mux12~19 (
// Equation(s):
// Mux122 = (temp_imemload_output_23 & ((\Mux12~16_combout  & (\Mux12~18_combout )) # (!\Mux12~16_combout  & ((\Mux12~11_combout ))))) # (!temp_imemload_output_23 & (((\Mux12~16_combout ))))

	.dataa(\Mux12~18_combout ),
	.datab(temp_imemload_output_23),
	.datac(\Mux12~16_combout ),
	.datad(\Mux12~11_combout ),
	.cin(gnd),
	.combout(Mux122),
	.cout());
// synopsys translate_off
defparam \Mux12~19 .lut_mask = 16'hBCB0;
defparam \Mux12~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N2
cycloneive_lcell_comb \Mux13~9 (
// Equation(s):
// Mux131 = (\Mux13~6_combout  & ((\Mux13~8_combout ) # ((!temp_imemload_output_21)))) # (!\Mux13~6_combout  & (((temp_imemload_output_21 & \Mux13~1_combout ))))

	.dataa(\Mux13~6_combout ),
	.datab(\Mux13~8_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux13~1_combout ),
	.cin(gnd),
	.combout(Mux131),
	.cout());
// synopsys translate_off
defparam \Mux13~9 .lut_mask = 16'hDA8A;
defparam \Mux13~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N14
cycloneive_lcell_comb \Mux13~19 (
// Equation(s):
// Mux132 = (temp_imemload_output_24 & ((\Mux13~16_combout  & (\Mux13~18_combout )) # (!\Mux13~16_combout  & ((\Mux13~11_combout ))))) # (!temp_imemload_output_24 & (((\Mux13~16_combout ))))

	.dataa(\Mux13~18_combout ),
	.datab(temp_imemload_output_24),
	.datac(\Mux13~11_combout ),
	.datad(\Mux13~16_combout ),
	.cin(gnd),
	.combout(Mux132),
	.cout());
// synopsys translate_off
defparam \Mux13~19 .lut_mask = 16'hBBC0;
defparam \Mux13~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N2
cycloneive_lcell_comb \Mux7~9 (
// Equation(s):
// Mux71 = (temp_imemload_output_21 & ((\Mux7~6_combout  & ((\Mux7~8_combout ))) # (!\Mux7~6_combout  & (\Mux7~1_combout )))) # (!temp_imemload_output_21 & (((\Mux7~6_combout ))))

	.dataa(\Mux7~1_combout ),
	.datab(\Mux7~8_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux7~6_combout ),
	.cin(gnd),
	.combout(Mux71),
	.cout());
// synopsys translate_off
defparam \Mux7~9 .lut_mask = 16'hCFA0;
defparam \Mux7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N24
cycloneive_lcell_comb \Mux7~19 (
// Equation(s):
// Mux72 = (\Mux7~16_combout  & ((\Mux7~18_combout ) # ((!temp_imemload_output_24)))) # (!\Mux7~16_combout  & (((\Mux7~11_combout  & temp_imemload_output_24))))

	.dataa(\Mux7~18_combout ),
	.datab(\Mux7~11_combout ),
	.datac(\Mux7~16_combout ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(Mux72),
	.cout());
// synopsys translate_off
defparam \Mux7~19 .lut_mask = 16'hACF0;
defparam \Mux7~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N24
cycloneive_lcell_comb \Mux8~9 (
// Equation(s):
// Mux81 = (\Mux8~6_combout  & (((\Mux8~8_combout ) # (!temp_imemload_output_21)))) # (!\Mux8~6_combout  & (\Mux8~1_combout  & (temp_imemload_output_21)))

	.dataa(\Mux8~6_combout ),
	.datab(\Mux8~1_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux8~8_combout ),
	.cin(gnd),
	.combout(Mux81),
	.cout());
// synopsys translate_off
defparam \Mux8~9 .lut_mask = 16'hEA4A;
defparam \Mux8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N12
cycloneive_lcell_comb \Mux8~19 (
// Equation(s):
// Mux82 = (\Mux8~16_combout  & (((\Mux8~18_combout ) # (!temp_imemload_output_23)))) # (!\Mux8~16_combout  & (\Mux8~11_combout  & (temp_imemload_output_23)))

	.dataa(\Mux8~11_combout ),
	.datab(\Mux8~16_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux8~18_combout ),
	.cin(gnd),
	.combout(Mux82),
	.cout());
// synopsys translate_off
defparam \Mux8~19 .lut_mask = 16'hEC2C;
defparam \Mux8~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N22
cycloneive_lcell_comb \Mux9~9 (
// Equation(s):
// Mux91 = (temp_imemload_output_21 & ((\Mux9~6_combout  & (\Mux9~8_combout )) # (!\Mux9~6_combout  & ((\Mux9~1_combout ))))) # (!temp_imemload_output_21 & (((\Mux9~6_combout ))))

	.dataa(\Mux9~8_combout ),
	.datab(\Mux9~1_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux9~6_combout ),
	.cin(gnd),
	.combout(Mux91),
	.cout());
// synopsys translate_off
defparam \Mux9~9 .lut_mask = 16'hAFC0;
defparam \Mux9~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N20
cycloneive_lcell_comb \Mux9~19 (
// Equation(s):
// Mux92 = (\Mux9~16_combout  & (((\Mux9~18_combout ) # (!temp_imemload_output_24)))) # (!\Mux9~16_combout  & (\Mux9~11_combout  & ((temp_imemload_output_24))))

	.dataa(\Mux9~11_combout ),
	.datab(\Mux9~18_combout ),
	.datac(\Mux9~16_combout ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(Mux92),
	.cout());
// synopsys translate_off
defparam \Mux9~19 .lut_mask = 16'hCAF0;
defparam \Mux9~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N18
cycloneive_lcell_comb \Mux10~9 (
// Equation(s):
// Mux101 = (\Mux10~6_combout  & (((\Mux10~8_combout ) # (!temp_imemload_output_21)))) # (!\Mux10~6_combout  & (\Mux10~1_combout  & ((temp_imemload_output_21))))

	.dataa(\Mux10~6_combout ),
	.datab(\Mux10~1_combout ),
	.datac(\Mux10~8_combout ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(Mux101),
	.cout());
// synopsys translate_off
defparam \Mux10~9 .lut_mask = 16'hE4AA;
defparam \Mux10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N2
cycloneive_lcell_comb \Mux10~19 (
// Equation(s):
// Mux102 = (\Mux10~16_combout  & ((\Mux10~18_combout ) # ((!temp_imemload_output_23)))) # (!\Mux10~16_combout  & (((temp_imemload_output_23 & \Mux10~11_combout ))))

	.dataa(\Mux10~16_combout ),
	.datab(\Mux10~18_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux10~11_combout ),
	.cin(gnd),
	.combout(Mux102),
	.cout());
// synopsys translate_off
defparam \Mux10~19 .lut_mask = 16'hDA8A;
defparam \Mux10~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N18
cycloneive_lcell_comb \Mux48~9 (
// Equation(s):
// Mux48 = (\Mux48~6_combout  & ((\Mux48~8_combout ) # ((!temp_imemload_output_16)))) # (!\Mux48~6_combout  & (((\Mux48~1_combout  & temp_imemload_output_16))))

	.dataa(\Mux48~6_combout ),
	.datab(\Mux48~8_combout ),
	.datac(\Mux48~1_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(Mux48),
	.cout());
// synopsys translate_off
defparam \Mux48~9 .lut_mask = 16'hD8AA;
defparam \Mux48~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N26
cycloneive_lcell_comb \Mux48~19 (
// Equation(s):
// Mux481 = (\Mux48~16_combout  & ((\Mux48~18_combout ) # ((!temp_imemload_output_19)))) # (!\Mux48~16_combout  & (((temp_imemload_output_19 & \Mux48~11_combout ))))

	.dataa(\Mux48~18_combout ),
	.datab(\Mux48~16_combout ),
	.datac(temp_imemload_output_19),
	.datad(\Mux48~11_combout ),
	.cin(gnd),
	.combout(Mux481),
	.cout());
// synopsys translate_off
defparam \Mux48~19 .lut_mask = 16'hBC8C;
defparam \Mux48~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N18
cycloneive_lcell_comb \Mux51~9 (
// Equation(s):
// Mux511 = (\Mux51~6_combout  & ((\Mux51~8_combout ) # ((!temp_imemload_output_16)))) # (!\Mux51~6_combout  & (((\Mux51~1_combout  & temp_imemload_output_16))))

	.dataa(\Mux51~8_combout ),
	.datab(\Mux51~1_combout ),
	.datac(\Mux51~6_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(Mux511),
	.cout());
// synopsys translate_off
defparam \Mux51~9 .lut_mask = 16'hACF0;
defparam \Mux51~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N0
cycloneive_lcell_comb \Mux51~19 (
// Equation(s):
// Mux512 = (temp_imemload_output_18 & ((\Mux51~16_combout  & (\Mux51~18_combout )) # (!\Mux51~16_combout  & ((\Mux51~11_combout ))))) # (!temp_imemload_output_18 & (\Mux51~16_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux51~16_combout ),
	.datac(\Mux51~18_combout ),
	.datad(\Mux51~11_combout ),
	.cin(gnd),
	.combout(Mux512),
	.cout());
// synopsys translate_off
defparam \Mux51~19 .lut_mask = 16'hE6C4;
defparam \Mux51~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N0
cycloneive_lcell_comb \Mux36~9 (
// Equation(s):
// Mux36 = (\Mux36~6_combout  & (((\Mux36~8_combout ) # (!temp_imemload_output_16)))) # (!\Mux36~6_combout  & (\Mux36~1_combout  & ((temp_imemload_output_16))))

	.dataa(\Mux36~6_combout ),
	.datab(\Mux36~1_combout ),
	.datac(\Mux36~8_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(Mux36),
	.cout());
// synopsys translate_off
defparam \Mux36~9 .lut_mask = 16'hE4AA;
defparam \Mux36~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N2
cycloneive_lcell_comb \Mux36~19 (
// Equation(s):
// Mux361 = (temp_imemload_output_18 & ((\Mux36~16_combout  & (\Mux36~18_combout )) # (!\Mux36~16_combout  & ((\Mux36~11_combout ))))) # (!temp_imemload_output_18 & (((\Mux36~16_combout ))))

	.dataa(\Mux36~18_combout ),
	.datab(\Mux36~11_combout ),
	.datac(temp_imemload_output_18),
	.datad(\Mux36~16_combout ),
	.cin(gnd),
	.combout(Mux361),
	.cout());
// synopsys translate_off
defparam \Mux36~19 .lut_mask = 16'hAFC0;
defparam \Mux36~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N20
cycloneive_lcell_comb \Mux45~9 (
// Equation(s):
// Mux45 = (temp_imemload_output_16 & ((\Mux45~6_combout  & (\Mux45~8_combout )) # (!\Mux45~6_combout  & ((\Mux45~1_combout ))))) # (!temp_imemload_output_16 & (((\Mux45~6_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux45~8_combout ),
	.datac(\Mux45~1_combout ),
	.datad(\Mux45~6_combout ),
	.cin(gnd),
	.combout(Mux45),
	.cout());
// synopsys translate_off
defparam \Mux45~9 .lut_mask = 16'hDDA0;
defparam \Mux45~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N14
cycloneive_lcell_comb \Mux45~19 (
// Equation(s):
// Mux451 = (\Mux45~16_combout  & (((\Mux45~18_combout )) # (!temp_imemload_output_18))) # (!\Mux45~16_combout  & (temp_imemload_output_18 & (\Mux45~11_combout )))

	.dataa(\Mux45~16_combout ),
	.datab(temp_imemload_output_18),
	.datac(\Mux45~11_combout ),
	.datad(\Mux45~18_combout ),
	.cin(gnd),
	.combout(Mux451),
	.cout());
// synopsys translate_off
defparam \Mux45~19 .lut_mask = 16'hEA62;
defparam \Mux45~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N30
cycloneive_lcell_comb \Mux46~9 (
// Equation(s):
// Mux46 = (temp_imemload_output_16 & ((\Mux46~6_combout  & (\Mux46~8_combout )) # (!\Mux46~6_combout  & ((\Mux46~1_combout ))))) # (!temp_imemload_output_16 & (((\Mux46~6_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux46~8_combout ),
	.datac(\Mux46~1_combout ),
	.datad(\Mux46~6_combout ),
	.cin(gnd),
	.combout(Mux46),
	.cout());
// synopsys translate_off
defparam \Mux46~9 .lut_mask = 16'hDDA0;
defparam \Mux46~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N8
cycloneive_lcell_comb \Mux46~19 (
// Equation(s):
// Mux461 = (temp_imemload_output_19 & ((\Mux46~16_combout  & (\Mux46~18_combout )) # (!\Mux46~16_combout  & ((\Mux46~11_combout ))))) # (!temp_imemload_output_19 & (((\Mux46~16_combout ))))

	.dataa(\Mux46~18_combout ),
	.datab(temp_imemload_output_19),
	.datac(\Mux46~16_combout ),
	.datad(\Mux46~11_combout ),
	.cin(gnd),
	.combout(Mux461),
	.cout());
// synopsys translate_off
defparam \Mux46~19 .lut_mask = 16'hBCB0;
defparam \Mux46~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N22
cycloneive_lcell_comb \Mux47~9 (
// Equation(s):
// Mux47 = (temp_imemload_output_16 & ((\Mux47~6_combout  & ((\Mux47~8_combout ))) # (!\Mux47~6_combout  & (\Mux47~1_combout )))) # (!temp_imemload_output_16 & (((\Mux47~6_combout ))))

	.dataa(\Mux47~1_combout ),
	.datab(\Mux47~8_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux47~6_combout ),
	.cin(gnd),
	.combout(Mux47),
	.cout());
// synopsys translate_off
defparam \Mux47~9 .lut_mask = 16'hCFA0;
defparam \Mux47~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N18
cycloneive_lcell_comb \Mux47~19 (
// Equation(s):
// Mux471 = (temp_imemload_output_18 & ((\Mux47~16_combout  & ((\Mux47~18_combout ))) # (!\Mux47~16_combout  & (\Mux47~11_combout )))) # (!temp_imemload_output_18 & (\Mux47~16_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux47~16_combout ),
	.datac(\Mux47~11_combout ),
	.datad(\Mux47~18_combout ),
	.cin(gnd),
	.combout(Mux471),
	.cout());
// synopsys translate_off
defparam \Mux47~19 .lut_mask = 16'hEC64;
defparam \Mux47~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N30
cycloneive_lcell_comb \Mux32~9 (
// Equation(s):
// Mux321 = (\Mux32~6_combout  & (((\Mux32~8_combout ) # (!temp_imemload_output_16)))) # (!\Mux32~6_combout  & (\Mux32~1_combout  & ((temp_imemload_output_16))))

	.dataa(\Mux32~1_combout ),
	.datab(\Mux32~8_combout ),
	.datac(\Mux32~6_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(Mux321),
	.cout());
// synopsys translate_off
defparam \Mux32~9 .lut_mask = 16'hCAF0;
defparam \Mux32~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N28
cycloneive_lcell_comb \Mux32~19 (
// Equation(s):
// Mux322 = (\Mux32~16_combout  & (((\Mux32~18_combout ) # (!temp_imemload_output_19)))) # (!\Mux32~16_combout  & (\Mux32~11_combout  & ((temp_imemload_output_19))))

	.dataa(\Mux32~11_combout ),
	.datab(\Mux32~18_combout ),
	.datac(\Mux32~16_combout ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(Mux322),
	.cout());
// synopsys translate_off
defparam \Mux32~19 .lut_mask = 16'hCAF0;
defparam \Mux32~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N6
cycloneive_lcell_comb \Mux33~9 (
// Equation(s):
// Mux331 = (\Mux33~6_combout  & (((\Mux33~8_combout ) # (!temp_imemload_output_16)))) # (!\Mux33~6_combout  & (\Mux33~1_combout  & (temp_imemload_output_16)))

	.dataa(\Mux33~1_combout ),
	.datab(\Mux33~6_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux33~8_combout ),
	.cin(gnd),
	.combout(Mux331),
	.cout());
// synopsys translate_off
defparam \Mux33~9 .lut_mask = 16'hEC2C;
defparam \Mux33~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N10
cycloneive_lcell_comb \Mux33~19 (
// Equation(s):
// Mux332 = (temp_imemload_output_18 & ((\Mux33~16_combout  & ((\Mux33~18_combout ))) # (!\Mux33~16_combout  & (\Mux33~11_combout )))) # (!temp_imemload_output_18 & (((\Mux33~16_combout ))))

	.dataa(\Mux33~11_combout ),
	.datab(\Mux33~18_combout ),
	.datac(temp_imemload_output_18),
	.datad(\Mux33~16_combout ),
	.cin(gnd),
	.combout(Mux332),
	.cout());
// synopsys translate_off
defparam \Mux33~19 .lut_mask = 16'hCFA0;
defparam \Mux33~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N16
cycloneive_lcell_comb \Mux34~9 (
// Equation(s):
// Mux34 = (\Mux34~6_combout  & ((\Mux34~8_combout ) # ((!temp_imemload_output_16)))) # (!\Mux34~6_combout  & (((temp_imemload_output_16 & \Mux34~1_combout ))))

	.dataa(\Mux34~8_combout ),
	.datab(\Mux34~6_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux34~1_combout ),
	.cin(gnd),
	.combout(Mux34),
	.cout());
// synopsys translate_off
defparam \Mux34~9 .lut_mask = 16'hBC8C;
defparam \Mux34~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N2
cycloneive_lcell_comb \Mux34~19 (
// Equation(s):
// Mux341 = (temp_imemload_output_19 & ((\Mux34~16_combout  & ((\Mux34~18_combout ))) # (!\Mux34~16_combout  & (\Mux34~11_combout )))) # (!temp_imemload_output_19 & (((\Mux34~16_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\Mux34~11_combout ),
	.datac(\Mux34~16_combout ),
	.datad(\Mux34~18_combout ),
	.cin(gnd),
	.combout(Mux341),
	.cout());
// synopsys translate_off
defparam \Mux34~19 .lut_mask = 16'hF858;
defparam \Mux34~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N4
cycloneive_lcell_comb \Mux35~9 (
// Equation(s):
// Mux35 = (temp_imemload_output_16 & ((\Mux35~6_combout  & (\Mux35~8_combout )) # (!\Mux35~6_combout  & ((\Mux35~1_combout ))))) # (!temp_imemload_output_16 & (((\Mux35~6_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux35~8_combout ),
	.datac(\Mux35~6_combout ),
	.datad(\Mux35~1_combout ),
	.cin(gnd),
	.combout(Mux35),
	.cout());
// synopsys translate_off
defparam \Mux35~9 .lut_mask = 16'hDAD0;
defparam \Mux35~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N4
cycloneive_lcell_comb \Mux35~19 (
// Equation(s):
// Mux351 = (temp_imemload_output_18 & ((\Mux35~16_combout  & ((\Mux35~18_combout ))) # (!\Mux35~16_combout  & (\Mux35~11_combout )))) # (!temp_imemload_output_18 & (((\Mux35~16_combout ))))

	.dataa(\Mux35~11_combout ),
	.datab(temp_imemload_output_18),
	.datac(\Mux35~16_combout ),
	.datad(\Mux35~18_combout ),
	.cin(gnd),
	.combout(Mux351),
	.cout());
// synopsys translate_off
defparam \Mux35~19 .lut_mask = 16'hF838;
defparam \Mux35~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N16
cycloneive_lcell_comb \Mux37~9 (
// Equation(s):
// Mux37 = (temp_imemload_output_16 & ((\Mux37~6_combout  & ((\Mux37~8_combout ))) # (!\Mux37~6_combout  & (\Mux37~1_combout )))) # (!temp_imemload_output_16 & (((\Mux37~6_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux37~1_combout ),
	.datac(\Mux37~6_combout ),
	.datad(\Mux37~8_combout ),
	.cin(gnd),
	.combout(Mux37),
	.cout());
// synopsys translate_off
defparam \Mux37~9 .lut_mask = 16'hF858;
defparam \Mux37~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N16
cycloneive_lcell_comb \Mux37~19 (
// Equation(s):
// Mux371 = (\Mux37~16_combout  & (((\Mux37~18_combout ) # (!temp_imemload_output_18)))) # (!\Mux37~16_combout  & (\Mux37~11_combout  & ((temp_imemload_output_18))))

	.dataa(\Mux37~16_combout ),
	.datab(\Mux37~11_combout ),
	.datac(\Mux37~18_combout ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(Mux371),
	.cout());
// synopsys translate_off
defparam \Mux37~19 .lut_mask = 16'hE4AA;
defparam \Mux37~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N0
cycloneive_lcell_comb \Mux38~9 (
// Equation(s):
// Mux38 = (temp_imemload_output_16 & ((\Mux38~6_combout  & (\Mux38~8_combout )) # (!\Mux38~6_combout  & ((\Mux38~1_combout ))))) # (!temp_imemload_output_16 & (((\Mux38~6_combout ))))

	.dataa(\Mux38~8_combout ),
	.datab(temp_imemload_output_16),
	.datac(\Mux38~1_combout ),
	.datad(\Mux38~6_combout ),
	.cin(gnd),
	.combout(Mux38),
	.cout());
// synopsys translate_off
defparam \Mux38~9 .lut_mask = 16'hBBC0;
defparam \Mux38~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N24
cycloneive_lcell_comb \Mux38~19 (
// Equation(s):
// Mux381 = (\Mux38~16_combout  & ((\Mux38~18_combout ) # ((!temp_imemload_output_19)))) # (!\Mux38~16_combout  & (((temp_imemload_output_19 & \Mux38~11_combout ))))

	.dataa(\Mux38~16_combout ),
	.datab(\Mux38~18_combout ),
	.datac(temp_imemload_output_19),
	.datad(\Mux38~11_combout ),
	.cin(gnd),
	.combout(Mux381),
	.cout());
// synopsys translate_off
defparam \Mux38~19 .lut_mask = 16'hDA8A;
defparam \Mux38~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N6
cycloneive_lcell_comb \Mux39~9 (
// Equation(s):
// Mux39 = (\Mux39~6_combout  & (((\Mux39~8_combout ) # (!temp_imemload_output_16)))) # (!\Mux39~6_combout  & (\Mux39~1_combout  & ((temp_imemload_output_16))))

	.dataa(\Mux39~6_combout ),
	.datab(\Mux39~1_combout ),
	.datac(\Mux39~8_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(Mux39),
	.cout());
// synopsys translate_off
defparam \Mux39~9 .lut_mask = 16'hE4AA;
defparam \Mux39~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N28
cycloneive_lcell_comb \Mux39~19 (
// Equation(s):
// Mux391 = (temp_imemload_output_18 & ((\Mux39~16_combout  & ((\Mux39~18_combout ))) # (!\Mux39~16_combout  & (\Mux39~11_combout )))) # (!temp_imemload_output_18 & (((\Mux39~16_combout ))))

	.dataa(\Mux39~11_combout ),
	.datab(temp_imemload_output_18),
	.datac(\Mux39~18_combout ),
	.datad(\Mux39~16_combout ),
	.cin(gnd),
	.combout(Mux391),
	.cout());
// synopsys translate_off
defparam \Mux39~19 .lut_mask = 16'hF388;
defparam \Mux39~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N28
cycloneive_lcell_comb \Mux40~9 (
// Equation(s):
// Mux40 = (\Mux40~6_combout  & ((\Mux40~8_combout ) # ((!temp_imemload_output_16)))) # (!\Mux40~6_combout  & (((temp_imemload_output_16 & \Mux40~1_combout ))))

	.dataa(\Mux40~6_combout ),
	.datab(\Mux40~8_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux40~1_combout ),
	.cin(gnd),
	.combout(Mux40),
	.cout());
// synopsys translate_off
defparam \Mux40~9 .lut_mask = 16'hDA8A;
defparam \Mux40~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N28
cycloneive_lcell_comb \Mux40~19 (
// Equation(s):
// Mux401 = (temp_imemload_output_19 & ((\Mux40~16_combout  & (\Mux40~18_combout )) # (!\Mux40~16_combout  & ((\Mux40~11_combout ))))) # (!temp_imemload_output_19 & (((\Mux40~16_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\Mux40~18_combout ),
	.datac(\Mux40~16_combout ),
	.datad(\Mux40~11_combout ),
	.cin(gnd),
	.combout(Mux401),
	.cout());
// synopsys translate_off
defparam \Mux40~19 .lut_mask = 16'hDAD0;
defparam \Mux40~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N24
cycloneive_lcell_comb \Mux41~9 (
// Equation(s):
// Mux411 = (temp_imemload_output_16 & ((\Mux41~6_combout  & (\Mux41~8_combout )) # (!\Mux41~6_combout  & ((\Mux41~1_combout ))))) # (!temp_imemload_output_16 & (((\Mux41~6_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux41~8_combout ),
	.datac(\Mux41~6_combout ),
	.datad(\Mux41~1_combout ),
	.cin(gnd),
	.combout(Mux411),
	.cout());
// synopsys translate_off
defparam \Mux41~9 .lut_mask = 16'hDAD0;
defparam \Mux41~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N6
cycloneive_lcell_comb \Mux41~19 (
// Equation(s):
// Mux412 = (temp_imemload_output_18 & ((\Mux41~16_combout  & (\Mux41~18_combout )) # (!\Mux41~16_combout  & ((\Mux41~11_combout ))))) # (!temp_imemload_output_18 & (((\Mux41~16_combout ))))

	.dataa(\Mux41~18_combout ),
	.datab(temp_imemload_output_18),
	.datac(\Mux41~11_combout ),
	.datad(\Mux41~16_combout ),
	.cin(gnd),
	.combout(Mux412),
	.cout());
// synopsys translate_off
defparam \Mux41~19 .lut_mask = 16'hBBC0;
defparam \Mux41~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N16
cycloneive_lcell_comb \Mux42~9 (
// Equation(s):
// Mux421 = (\Mux42~6_combout  & ((\Mux42~8_combout ) # ((!temp_imemload_output_16)))) # (!\Mux42~6_combout  & (((\Mux42~1_combout  & temp_imemload_output_16))))

	.dataa(\Mux42~8_combout ),
	.datab(\Mux42~6_combout ),
	.datac(\Mux42~1_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(Mux421),
	.cout());
// synopsys translate_off
defparam \Mux42~9 .lut_mask = 16'hB8CC;
defparam \Mux42~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N14
cycloneive_lcell_comb \Mux42~19 (
// Equation(s):
// Mux422 = (\Mux42~16_combout  & ((\Mux42~18_combout ) # ((!temp_imemload_output_19)))) # (!\Mux42~16_combout  & (((temp_imemload_output_19 & \Mux42~11_combout ))))

	.dataa(\Mux42~16_combout ),
	.datab(\Mux42~18_combout ),
	.datac(temp_imemload_output_19),
	.datad(\Mux42~11_combout ),
	.cin(gnd),
	.combout(Mux422),
	.cout());
// synopsys translate_off
defparam \Mux42~19 .lut_mask = 16'hDA8A;
defparam \Mux42~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N20
cycloneive_lcell_comb \Mux43~9 (
// Equation(s):
// Mux43 = (temp_imemload_output_16 & ((\Mux43~6_combout  & ((\Mux43~8_combout ))) # (!\Mux43~6_combout  & (\Mux43~1_combout )))) # (!temp_imemload_output_16 & (((\Mux43~6_combout ))))

	.dataa(\Mux43~1_combout ),
	.datab(temp_imemload_output_16),
	.datac(\Mux43~6_combout ),
	.datad(\Mux43~8_combout ),
	.cin(gnd),
	.combout(Mux43),
	.cout());
// synopsys translate_off
defparam \Mux43~9 .lut_mask = 16'hF838;
defparam \Mux43~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N14
cycloneive_lcell_comb \Mux43~19 (
// Equation(s):
// Mux431 = (temp_imemload_output_18 & ((\Mux43~16_combout  & ((\Mux43~18_combout ))) # (!\Mux43~16_combout  & (\Mux43~11_combout )))) # (!temp_imemload_output_18 & (((\Mux43~16_combout ))))

	.dataa(\Mux43~11_combout ),
	.datab(temp_imemload_output_18),
	.datac(\Mux43~16_combout ),
	.datad(\Mux43~18_combout ),
	.cin(gnd),
	.combout(Mux431),
	.cout());
// synopsys translate_off
defparam \Mux43~19 .lut_mask = 16'hF838;
defparam \Mux43~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N2
cycloneive_lcell_comb \Mux44~9 (
// Equation(s):
// Mux44 = (temp_imemload_output_16 & ((\Mux44~6_combout  & (\Mux44~8_combout )) # (!\Mux44~6_combout  & ((\Mux44~1_combout ))))) # (!temp_imemload_output_16 & (((\Mux44~6_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux44~8_combout ),
	.datac(\Mux44~1_combout ),
	.datad(\Mux44~6_combout ),
	.cin(gnd),
	.combout(Mux44),
	.cout());
// synopsys translate_off
defparam \Mux44~9 .lut_mask = 16'hDDA0;
defparam \Mux44~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N30
cycloneive_lcell_comb \Mux44~19 (
// Equation(s):
// Mux441 = (temp_imemload_output_19 & ((\Mux44~16_combout  & ((\Mux44~18_combout ))) # (!\Mux44~16_combout  & (\Mux44~11_combout )))) # (!temp_imemload_output_19 & (((\Mux44~16_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\Mux44~11_combout ),
	.datac(\Mux44~16_combout ),
	.datad(\Mux44~18_combout ),
	.cin(gnd),
	.combout(Mux441),
	.cout());
// synopsys translate_off
defparam \Mux44~19 .lut_mask = 16'hF858;
defparam \Mux44~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N10
cycloneive_lcell_comb \Mux53~9 (
// Equation(s):
// Mux53 = (\Mux53~6_combout  & ((\Mux53~8_combout ) # ((!temp_imemload_output_16)))) # (!\Mux53~6_combout  & (((temp_imemload_output_16 & \Mux53~1_combout ))))

	.dataa(\Mux53~6_combout ),
	.datab(\Mux53~8_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux53~1_combout ),
	.cin(gnd),
	.combout(Mux53),
	.cout());
// synopsys translate_off
defparam \Mux53~9 .lut_mask = 16'hDA8A;
defparam \Mux53~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N4
cycloneive_lcell_comb \Mux53~19 (
// Equation(s):
// Mux531 = (temp_imemload_output_19 & ((\Mux53~16_combout  & (\Mux53~18_combout )) # (!\Mux53~16_combout  & ((\Mux53~11_combout ))))) # (!temp_imemload_output_19 & (((\Mux53~16_combout ))))

	.dataa(\Mux53~18_combout ),
	.datab(\Mux53~11_combout ),
	.datac(temp_imemload_output_19),
	.datad(\Mux53~16_combout ),
	.cin(gnd),
	.combout(Mux531),
	.cout());
// synopsys translate_off
defparam \Mux53~19 .lut_mask = 16'hAFC0;
defparam \Mux53~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N20
cycloneive_lcell_comb \Mux49~9 (
// Equation(s):
// Mux49 = (temp_imemload_output_16 & ((\Mux49~6_combout  & (\Mux49~8_combout )) # (!\Mux49~6_combout  & ((\Mux49~1_combout ))))) # (!temp_imemload_output_16 & (((\Mux49~6_combout ))))

	.dataa(\Mux49~8_combout ),
	.datab(temp_imemload_output_16),
	.datac(\Mux49~1_combout ),
	.datad(\Mux49~6_combout ),
	.cin(gnd),
	.combout(Mux49),
	.cout());
// synopsys translate_off
defparam \Mux49~9 .lut_mask = 16'hBBC0;
defparam \Mux49~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N8
cycloneive_lcell_comb \Mux49~19 (
// Equation(s):
// Mux491 = (temp_imemload_output_18 & ((\Mux49~16_combout  & (\Mux49~18_combout )) # (!\Mux49~16_combout  & ((\Mux49~11_combout ))))) # (!temp_imemload_output_18 & (((\Mux49~16_combout ))))

	.dataa(\Mux49~18_combout ),
	.datab(temp_imemload_output_18),
	.datac(\Mux49~16_combout ),
	.datad(\Mux49~11_combout ),
	.cin(gnd),
	.combout(Mux491),
	.cout());
// synopsys translate_off
defparam \Mux49~19 .lut_mask = 16'hBCB0;
defparam \Mux49~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N4
cycloneive_lcell_comb \Mux54~9 (
// Equation(s):
// Mux54 = (\Mux54~6_combout  & ((\Mux54~8_combout ) # ((!temp_imemload_output_16)))) # (!\Mux54~6_combout  & (((\Mux54~1_combout  & temp_imemload_output_16))))

	.dataa(\Mux54~8_combout ),
	.datab(\Mux54~1_combout ),
	.datac(\Mux54~6_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(Mux54),
	.cout());
// synopsys translate_off
defparam \Mux54~9 .lut_mask = 16'hACF0;
defparam \Mux54~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N4
cycloneive_lcell_comb \Mux54~19 (
// Equation(s):
// Mux541 = (\Mux54~16_combout  & ((\Mux54~18_combout ) # ((!temp_imemload_output_19)))) # (!\Mux54~16_combout  & (((\Mux54~11_combout  & temp_imemload_output_19))))

	.dataa(\Mux54~18_combout ),
	.datab(\Mux54~16_combout ),
	.datac(\Mux54~11_combout ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(Mux541),
	.cout());
// synopsys translate_off
defparam \Mux54~19 .lut_mask = 16'hB8CC;
defparam \Mux54~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N0
cycloneive_lcell_comb \Mux55~9 (
// Equation(s):
// Mux55 = (temp_imemload_output_16 & ((\Mux55~6_combout  & (\Mux55~8_combout )) # (!\Mux55~6_combout  & ((\Mux55~1_combout ))))) # (!temp_imemload_output_16 & (((\Mux55~6_combout ))))

	.dataa(\Mux55~8_combout ),
	.datab(\Mux55~1_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux55~6_combout ),
	.cin(gnd),
	.combout(Mux55),
	.cout());
// synopsys translate_off
defparam \Mux55~9 .lut_mask = 16'hAFC0;
defparam \Mux55~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N24
cycloneive_lcell_comb \Mux55~19 (
// Equation(s):
// Mux551 = (temp_imemload_output_18 & ((\Mux55~16_combout  & (\Mux55~18_combout )) # (!\Mux55~16_combout  & ((\Mux55~11_combout ))))) # (!temp_imemload_output_18 & (((\Mux55~16_combout ))))

	.dataa(\Mux55~18_combout ),
	.datab(temp_imemload_output_18),
	.datac(\Mux55~11_combout ),
	.datad(\Mux55~16_combout ),
	.cin(gnd),
	.combout(Mux551),
	.cout());
// synopsys translate_off
defparam \Mux55~19 .lut_mask = 16'hBBC0;
defparam \Mux55~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N10
cycloneive_lcell_comb \Mux56~9 (
// Equation(s):
// Mux56 = (temp_imemload_output_16 & ((\Mux56~6_combout  & ((\Mux56~8_combout ))) # (!\Mux56~6_combout  & (\Mux56~1_combout )))) # (!temp_imemload_output_16 & (((\Mux56~6_combout ))))

	.dataa(\Mux56~1_combout ),
	.datab(\Mux56~8_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux56~6_combout ),
	.cin(gnd),
	.combout(Mux56),
	.cout());
// synopsys translate_off
defparam \Mux56~9 .lut_mask = 16'hCFA0;
defparam \Mux56~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N6
cycloneive_lcell_comb \Mux56~19 (
// Equation(s):
// Mux561 = (temp_imemload_output_19 & ((\Mux56~16_combout  & (\Mux56~18_combout )) # (!\Mux56~16_combout  & ((\Mux56~11_combout ))))) # (!temp_imemload_output_19 & (((\Mux56~16_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\Mux56~18_combout ),
	.datac(\Mux56~16_combout ),
	.datad(\Mux56~11_combout ),
	.cin(gnd),
	.combout(Mux561),
	.cout());
// synopsys translate_off
defparam \Mux56~19 .lut_mask = 16'hDAD0;
defparam \Mux56~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N2
cycloneive_lcell_comb \Mux57~9 (
// Equation(s):
// Mux57 = (temp_imemload_output_16 & ((\Mux57~6_combout  & (\Mux57~8_combout )) # (!\Mux57~6_combout  & ((\Mux57~1_combout ))))) # (!temp_imemload_output_16 & (((\Mux57~6_combout ))))

	.dataa(\Mux57~8_combout ),
	.datab(temp_imemload_output_16),
	.datac(\Mux57~6_combout ),
	.datad(\Mux57~1_combout ),
	.cin(gnd),
	.combout(Mux57),
	.cout());
// synopsys translate_off
defparam \Mux57~9 .lut_mask = 16'hBCB0;
defparam \Mux57~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N28
cycloneive_lcell_comb \Mux57~19 (
// Equation(s):
// Mux571 = (\Mux57~16_combout  & (((\Mux57~18_combout )) # (!temp_imemload_output_18))) # (!\Mux57~16_combout  & (temp_imemload_output_18 & (\Mux57~11_combout )))

	.dataa(\Mux57~16_combout ),
	.datab(temp_imemload_output_18),
	.datac(\Mux57~11_combout ),
	.datad(\Mux57~18_combout ),
	.cin(gnd),
	.combout(Mux571),
	.cout());
// synopsys translate_off
defparam \Mux57~19 .lut_mask = 16'hEA62;
defparam \Mux57~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N10
cycloneive_lcell_comb \Mux58~9 (
// Equation(s):
// Mux58 = (temp_imemload_output_16 & ((\Mux58~6_combout  & ((\Mux58~8_combout ))) # (!\Mux58~6_combout  & (\Mux58~1_combout )))) # (!temp_imemload_output_16 & (((\Mux58~6_combout ))))

	.dataa(\Mux58~1_combout ),
	.datab(temp_imemload_output_16),
	.datac(\Mux58~8_combout ),
	.datad(\Mux58~6_combout ),
	.cin(gnd),
	.combout(Mux58),
	.cout());
// synopsys translate_off
defparam \Mux58~9 .lut_mask = 16'hF388;
defparam \Mux58~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N4
cycloneive_lcell_comb \Mux58~19 (
// Equation(s):
// Mux581 = (temp_imemload_output_19 & ((\Mux58~16_combout  & (\Mux58~18_combout )) # (!\Mux58~16_combout  & ((\Mux58~11_combout ))))) # (!temp_imemload_output_19 & (((\Mux58~16_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\Mux58~18_combout ),
	.datac(\Mux58~11_combout ),
	.datad(\Mux58~16_combout ),
	.cin(gnd),
	.combout(Mux581),
	.cout());
// synopsys translate_off
defparam \Mux58~19 .lut_mask = 16'hDDA0;
defparam \Mux58~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N26
cycloneive_lcell_comb \Mux50~9 (
// Equation(s):
// Mux50 = (temp_imemload_output_16 & ((\Mux50~6_combout  & (\Mux50~8_combout )) # (!\Mux50~6_combout  & ((\Mux50~1_combout ))))) # (!temp_imemload_output_16 & (((\Mux50~6_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux50~8_combout ),
	.datac(\Mux50~6_combout ),
	.datad(\Mux50~1_combout ),
	.cin(gnd),
	.combout(Mux50),
	.cout());
// synopsys translate_off
defparam \Mux50~9 .lut_mask = 16'hDAD0;
defparam \Mux50~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N30
cycloneive_lcell_comb \Mux50~19 (
// Equation(s):
// Mux501 = (temp_imemload_output_19 & ((\Mux50~16_combout  & ((\Mux50~18_combout ))) # (!\Mux50~16_combout  & (\Mux50~11_combout )))) # (!temp_imemload_output_19 & (((\Mux50~16_combout ))))

	.dataa(\Mux50~11_combout ),
	.datab(temp_imemload_output_19),
	.datac(\Mux50~16_combout ),
	.datad(\Mux50~18_combout ),
	.cin(gnd),
	.combout(Mux501),
	.cout());
// synopsys translate_off
defparam \Mux50~19 .lut_mask = 16'hF838;
defparam \Mux50~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N20
cycloneive_lcell_comb \Mux52~9 (
// Equation(s):
// Mux521 = (\Mux52~6_combout  & ((\Mux52~8_combout ) # ((!temp_imemload_output_16)))) # (!\Mux52~6_combout  & (((\Mux52~1_combout  & temp_imemload_output_16))))

	.dataa(\Mux52~8_combout ),
	.datab(\Mux52~6_combout ),
	.datac(\Mux52~1_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(Mux521),
	.cout());
// synopsys translate_off
defparam \Mux52~9 .lut_mask = 16'hB8CC;
defparam \Mux52~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N22
cycloneive_lcell_comb \Mux52~19 (
// Equation(s):
// Mux522 = (\Mux52~16_combout  & ((\Mux52~18_combout ) # ((!temp_imemload_output_19)))) # (!\Mux52~16_combout  & (((\Mux52~11_combout  & temp_imemload_output_19))))

	.dataa(\Mux52~16_combout ),
	.datab(\Mux52~18_combout ),
	.datac(\Mux52~11_combout ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(Mux522),
	.cout());
// synopsys translate_off
defparam \Mux52~19 .lut_mask = 16'hD8AA;
defparam \Mux52~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N12
cycloneive_lcell_comb \storeregister[31][1]~feeder (
// Equation(s):
// \storeregister[31][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux30),
	.cin(gnd),
	.combout(\storeregister[31][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][1]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[31][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N8
cycloneive_lcell_comb \Decoder0~9 (
// Equation(s):
// \Decoder0~9_combout  = (temp_branchDest_01 & (temp_regwrite2 & temp_branchDest_41))

	.dataa(temp_branchDest_0),
	.datab(temp_regwrite),
	.datac(gnd),
	.datad(temp_branchDest_4),
	.cin(gnd),
	.combout(\Decoder0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~9 .lut_mask = 16'h8800;
defparam \Decoder0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N10
cycloneive_lcell_comb \Decoder0~27 (
// Equation(s):
// \Decoder0~27_combout  = (temp_branchDest_31 & (temp_branchDest_21 & (temp_branchDest_11 & \Decoder0~9_combout )))

	.dataa(temp_branchDest_3),
	.datab(temp_branchDest_2),
	.datac(temp_branchDest_1),
	.datad(\Decoder0~9_combout ),
	.cin(gnd),
	.combout(\Decoder0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~27 .lut_mask = 16'h8000;
defparam \Decoder0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N13
dffeas \storeregister[31][1] (
	.clk(!CLK),
	.d(\storeregister[31][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][1] .is_wysiwyg = "true";
defparam \storeregister[31][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N8
cycloneive_lcell_comb \storeregister[27][1]~feeder (
// Equation(s):
// \storeregister[27][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux30),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][1]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N8
cycloneive_lcell_comb \Decoder0~25 (
// Equation(s):
// \Decoder0~25_combout  = (temp_branchDest_11 & (\Decoder0~9_combout  & (!temp_branchDest_21 & temp_branchDest_31)))

	.dataa(temp_branchDest_1),
	.datab(\Decoder0~9_combout ),
	.datac(temp_branchDest_2),
	.datad(temp_branchDest_3),
	.cin(gnd),
	.combout(\Decoder0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~25 .lut_mask = 16'h0800;
defparam \Decoder0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N9
dffeas \storeregister[27][1] (
	.clk(!CLK),
	.d(\storeregister[27][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][1] .is_wysiwyg = "true";
defparam \storeregister[27][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N28
cycloneive_lcell_comb \storeregister[19][1]~feeder (
// Equation(s):
// \storeregister[19][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux30),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[19][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[19][1]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[19][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N8
cycloneive_lcell_comb \Decoder0~26 (
// Equation(s):
// \Decoder0~26_combout  = (!temp_branchDest_31 & (!temp_branchDest_21 & (temp_branchDest_11 & \Decoder0~9_combout )))

	.dataa(temp_branchDest_3),
	.datab(temp_branchDest_2),
	.datac(temp_branchDest_1),
	.datad(\Decoder0~9_combout ),
	.cin(gnd),
	.combout(\Decoder0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~26 .lut_mask = 16'h1000;
defparam \Decoder0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N29
dffeas \storeregister[19][1] (
	.clk(!CLK),
	.d(\storeregister[19][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][1] .is_wysiwyg = "true";
defparam \storeregister[19][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N18
cycloneive_lcell_comb \Mux62~7 (
// Equation(s):
// \Mux62~7_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\storeregister[27][1]~q )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & ((\storeregister[19][1]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[27][1]~q ),
	.datad(\storeregister[19][1]~q ),
	.cin(gnd),
	.combout(\Mux62~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~7 .lut_mask = 16'hB9A8;
defparam \Mux62~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N16
cycloneive_lcell_comb \storeregister[23][1]~feeder (
// Equation(s):
// \storeregister[23][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux30),
	.cin(gnd),
	.combout(\storeregister[23][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][1]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[23][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N24
cycloneive_lcell_comb \Decoder0~24 (
// Equation(s):
// \Decoder0~24_combout  = (temp_branchDest_21 & (\Decoder0~9_combout  & (!temp_branchDest_31 & temp_branchDest_11)))

	.dataa(temp_branchDest_2),
	.datab(\Decoder0~9_combout ),
	.datac(temp_branchDest_3),
	.datad(temp_branchDest_1),
	.cin(gnd),
	.combout(\Decoder0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~24 .lut_mask = 16'h0800;
defparam \Decoder0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N17
dffeas \storeregister[23][1] (
	.clk(!CLK),
	.d(\storeregister[23][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][1] .is_wysiwyg = "true";
defparam \storeregister[23][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N30
cycloneive_lcell_comb \Mux62~8 (
// Equation(s):
// \Mux62~8_combout  = (\Mux62~7_combout  & ((\storeregister[31][1]~q ) # ((!temp_imemload_output_18)))) # (!\Mux62~7_combout  & (((temp_imemload_output_18 & \storeregister[23][1]~q ))))

	.dataa(\storeregister[31][1]~q ),
	.datab(\Mux62~7_combout ),
	.datac(temp_imemload_output_18),
	.datad(\storeregister[23][1]~q ),
	.cin(gnd),
	.combout(\Mux62~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~8 .lut_mask = 16'hBC8C;
defparam \Mux62~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N8
cycloneive_lcell_comb \storeregister[17][1]~feeder (
// Equation(s):
// \storeregister[17][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux30),
	.cin(gnd),
	.combout(\storeregister[17][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[17][1]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[17][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N14
cycloneive_lcell_comb \Decoder0~44 (
// Equation(s):
// \Decoder0~44_combout  = (!temp_branchDest_31 & (!temp_branchDest_21 & (!temp_branchDest_11 & \Decoder0~9_combout )))

	.dataa(temp_branchDest_3),
	.datab(temp_branchDest_2),
	.datac(temp_branchDest_1),
	.datad(\Decoder0~9_combout ),
	.cin(gnd),
	.combout(\Decoder0~44_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~44 .lut_mask = 16'h0100;
defparam \Decoder0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N9
dffeas \storeregister[17][1] (
	.clk(!CLK),
	.d(\storeregister[17][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][1] .is_wysiwyg = "true";
defparam \storeregister[17][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N26
cycloneive_lcell_comb \storeregister[25][1]~feeder (
// Equation(s):
// \storeregister[25][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux30),
	.cin(gnd),
	.combout(\storeregister[25][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[25][1]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[25][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N28
cycloneive_lcell_comb \Decoder0~10 (
// Equation(s):
// \Decoder0~10_combout  = (temp_branchDest_01 & (!temp_branchDest_11 & (temp_regwrite2 & temp_branchDest_31)))

	.dataa(temp_branchDest_0),
	.datab(temp_branchDest_1),
	.datac(temp_regwrite),
	.datad(temp_branchDest_3),
	.cin(gnd),
	.combout(\Decoder0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~10 .lut_mask = 16'h2000;
defparam \Decoder0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N2
cycloneive_lcell_comb \Decoder0~11 (
// Equation(s):
// \Decoder0~11_combout  = (!temp_branchDest_21 & (\Decoder0~10_combout  & temp_branchDest_41))

	.dataa(gnd),
	.datab(temp_branchDest_2),
	.datac(\Decoder0~10_combout ),
	.datad(temp_branchDest_4),
	.cin(gnd),
	.combout(\Decoder0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~11 .lut_mask = 16'h3000;
defparam \Decoder0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N27
dffeas \storeregister[25][1] (
	.clk(!CLK),
	.d(\storeregister[25][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][1] .is_wysiwyg = "true";
defparam \storeregister[25][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N22
cycloneive_lcell_comb \Mux62~0 (
// Equation(s):
// \Mux62~0_combout  = (temp_imemload_output_19 & (((\storeregister[25][1]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[17][1]~q  & ((!temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[17][1]~q ),
	.datac(\storeregister[25][1]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~0 .lut_mask = 16'hAAE4;
defparam \Mux62~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N0
cycloneive_lcell_comb \Decoder0~43 (
// Equation(s):
// \Decoder0~43_combout  = (!temp_branchDest_31 & (temp_branchDest_21 & (!temp_branchDest_11 & \Decoder0~9_combout )))

	.dataa(temp_branchDest_3),
	.datab(temp_branchDest_2),
	.datac(temp_branchDest_1),
	.datad(\Decoder0~9_combout ),
	.cin(gnd),
	.combout(\Decoder0~43_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~43 .lut_mask = 16'h0400;
defparam \Decoder0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N23
dffeas \storeregister[21][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][1] .is_wysiwyg = "true";
defparam \storeregister[21][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N8
cycloneive_lcell_comb \storeregister[29][1]~feeder (
// Equation(s):
// \storeregister[29][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux30),
	.cin(gnd),
	.combout(\storeregister[29][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][1]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[29][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N12
cycloneive_lcell_comb \Decoder0~12 (
// Equation(s):
// \Decoder0~12_combout  = (temp_branchDest_21 & (temp_branchDest_41 & \Decoder0~10_combout ))

	.dataa(temp_branchDest_2),
	.datab(gnd),
	.datac(temp_branchDest_4),
	.datad(\Decoder0~10_combout ),
	.cin(gnd),
	.combout(\Decoder0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~12 .lut_mask = 16'hA000;
defparam \Decoder0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N9
dffeas \storeregister[29][1] (
	.clk(!CLK),
	.d(\storeregister[29][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][1] .is_wysiwyg = "true";
defparam \storeregister[29][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N10
cycloneive_lcell_comb \Mux62~1 (
// Equation(s):
// \Mux62~1_combout  = (temp_imemload_output_18 & ((\Mux62~0_combout  & ((\storeregister[29][1]~q ))) # (!\Mux62~0_combout  & (\storeregister[21][1]~q )))) # (!temp_imemload_output_18 & (\Mux62~0_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux62~0_combout ),
	.datac(\storeregister[21][1]~q ),
	.datad(\storeregister[29][1]~q ),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~1 .lut_mask = 16'hEC64;
defparam \Mux62~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N28
cycloneive_lcell_comb \storeregister[26][1]~feeder (
// Equation(s):
// \storeregister[26][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux30),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[26][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[26][1]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[26][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N20
cycloneive_lcell_comb \Decoder0~14 (
// Equation(s):
// \Decoder0~14_combout  = (\Decoder0~13_combout  & (temp_branchDest_41 & (temp_branchDest_31 & !temp_branchDest_21)))

	.dataa(\Decoder0~13_combout ),
	.datab(temp_branchDest_4),
	.datac(temp_branchDest_3),
	.datad(temp_branchDest_2),
	.cin(gnd),
	.combout(\Decoder0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~14 .lut_mask = 16'h0080;
defparam \Decoder0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N29
dffeas \storeregister[26][1] (
	.clk(!CLK),
	.d(\storeregister[26][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][1] .is_wysiwyg = "true";
defparam \storeregister[26][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N4
cycloneive_lcell_comb \storeregister[30][1]~feeder (
// Equation(s):
// \storeregister[30][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux30),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[30][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][1]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[30][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N14
cycloneive_lcell_comb \Decoder0~17 (
// Equation(s):
// \Decoder0~17_combout  = (\Decoder0~13_combout  & (temp_branchDest_41 & (temp_branchDest_31 & temp_branchDest_21)))

	.dataa(\Decoder0~13_combout ),
	.datab(temp_branchDest_4),
	.datac(temp_branchDest_3),
	.datad(temp_branchDest_2),
	.cin(gnd),
	.combout(\Decoder0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~17 .lut_mask = 16'h8000;
defparam \Decoder0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N5
dffeas \storeregister[30][1] (
	.clk(!CLK),
	.d(\storeregister[30][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][1] .is_wysiwyg = "true";
defparam \storeregister[30][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N24
cycloneive_lcell_comb \Mux62~3 (
// Equation(s):
// \Mux62~3_combout  = (\Mux62~2_combout  & (((\storeregister[30][1]~q ) # (!temp_imemload_output_19)))) # (!\Mux62~2_combout  & (\storeregister[26][1]~q  & ((temp_imemload_output_19))))

	.dataa(\Mux62~2_combout ),
	.datab(\storeregister[26][1]~q ),
	.datac(\storeregister[30][1]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux62~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~3 .lut_mask = 16'hE4AA;
defparam \Mux62~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N12
cycloneive_lcell_comb \Decoder0~8 (
// Equation(s):
// \Decoder0~8_combout  = (!temp_branchDest_11 & !temp_branchDest_31)

	.dataa(gnd),
	.datab(temp_branchDest_1),
	.datac(gnd),
	.datad(temp_branchDest_3),
	.cin(gnd),
	.combout(\Decoder0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~8 .lut_mask = 16'h0033;
defparam \Decoder0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N22
cycloneive_lcell_comb \Decoder0~21 (
// Equation(s):
// \Decoder0~21_combout  = (\Decoder0~20_combout  & (temp_branchDest_41 & (\Decoder0~8_combout  & temp_branchDest_21)))

	.dataa(\Decoder0~20_combout ),
	.datab(temp_branchDest_4),
	.datac(\Decoder0~8_combout ),
	.datad(temp_branchDest_2),
	.cin(gnd),
	.combout(\Decoder0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~21 .lut_mask = 16'h8000;
defparam \Decoder0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N21
dffeas \storeregister[20][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][1] .is_wysiwyg = "true";
defparam \storeregister[20][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N4
cycloneive_lcell_comb \Decoder0~22 (
// Equation(s):
// \Decoder0~22_combout  = (\Decoder0~20_combout  & (temp_branchDest_41 & (\Decoder0~8_combout  & !temp_branchDest_21)))

	.dataa(\Decoder0~20_combout ),
	.datab(temp_branchDest_4),
	.datac(\Decoder0~8_combout ),
	.datad(temp_branchDest_2),
	.cin(gnd),
	.combout(\Decoder0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~22 .lut_mask = 16'h0080;
defparam \Decoder0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N3
dffeas \storeregister[16][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][1] .is_wysiwyg = "true";
defparam \storeregister[16][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N20
cycloneive_lcell_comb \Mux62~4 (
// Equation(s):
// \Mux62~4_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\storeregister[20][1]~q )) # (!temp_imemload_output_18 & ((\storeregister[16][1]~q )))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[20][1]~q ),
	.datad(\storeregister[16][1]~q ),
	.cin(gnd),
	.combout(\Mux62~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~4 .lut_mask = 16'hD9C8;
defparam \Mux62~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N20
cycloneive_lcell_comb \storeregister[24][1]~feeder (
// Equation(s):
// \storeregister[24][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux30),
	.cin(gnd),
	.combout(\storeregister[24][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][1]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[24][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N12
cycloneive_lcell_comb \Decoder0~19 (
// Equation(s):
// \Decoder0~19_combout  = (\Decoder0~18_combout  & (!temp_branchDest_21 & temp_branchDest_41))

	.dataa(\Decoder0~18_combout ),
	.datab(temp_branchDest_2),
	.datac(gnd),
	.datad(temp_branchDest_4),
	.cin(gnd),
	.combout(\Decoder0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~19 .lut_mask = 16'h2200;
defparam \Decoder0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N21
dffeas \storeregister[24][1] (
	.clk(!CLK),
	.d(\storeregister[24][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][1] .is_wysiwyg = "true";
defparam \storeregister[24][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N24
cycloneive_lcell_comb \Mux62~5 (
// Equation(s):
// \Mux62~5_combout  = (\Mux62~4_combout  & ((\storeregister[28][1]~q ) # ((!temp_imemload_output_19)))) # (!\Mux62~4_combout  & (((temp_imemload_output_19 & \storeregister[24][1]~q ))))

	.dataa(\storeregister[28][1]~q ),
	.datab(\Mux62~4_combout ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[24][1]~q ),
	.cin(gnd),
	.combout(\Mux62~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~5 .lut_mask = 16'hBC8C;
defparam \Mux62~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N24
cycloneive_lcell_comb \Mux62~6 (
// Equation(s):
// \Mux62~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\Mux62~3_combout )) # (!temp_imemload_output_17 & ((\Mux62~5_combout )))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux62~3_combout ),
	.datac(temp_imemload_output_17),
	.datad(\Mux62~5_combout ),
	.cin(gnd),
	.combout(\Mux62~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~6 .lut_mask = 16'hE5E0;
defparam \Mux62~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N14
cycloneive_lcell_comb \Decoder0~30 (
// Equation(s):
// \Decoder0~30_combout  = (temp_branchDest_01 & (temp_regwrite2 & !temp_branchDest_41))

	.dataa(temp_branchDest_0),
	.datab(temp_regwrite),
	.datac(gnd),
	.datad(temp_branchDest_4),
	.cin(gnd),
	.combout(\Decoder0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~30 .lut_mask = 16'h0088;
defparam \Decoder0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N0
cycloneive_lcell_comb \Decoder0~45 (
// Equation(s):
// \Decoder0~45_combout  = (!temp_branchDest_11 & (!temp_branchDest_31 & (temp_branchDest_21 & \Decoder0~30_combout )))

	.dataa(temp_branchDest_1),
	.datab(temp_branchDest_3),
	.datac(temp_branchDest_2),
	.datad(\Decoder0~30_combout ),
	.cin(gnd),
	.combout(\Decoder0~45_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~45 .lut_mask = 16'h1000;
defparam \Decoder0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y42_N5
dffeas \storeregister[5][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][1] .is_wysiwyg = "true";
defparam \storeregister[5][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N4
cycloneive_lcell_comb \Mux62~10 (
// Equation(s):
// \Mux62~10_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[5][1]~q ))) # (!temp_imemload_output_16 & (\storeregister[4][1]~q ))))

	.dataa(\storeregister[4][1]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][1]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux62~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~10 .lut_mask = 16'hFC22;
defparam \Mux62~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N28
cycloneive_lcell_comb \storeregister[7][1]~feeder (
// Equation(s):
// \storeregister[7][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux30),
	.cin(gnd),
	.combout(\storeregister[7][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[7][1]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[7][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N30
cycloneive_lcell_comb \Decoder0~32 (
// Equation(s):
// \Decoder0~32_combout  = (temp_branchDest_11 & (!temp_branchDest_31 & (temp_branchDest_21 & \Decoder0~30_combout )))

	.dataa(temp_branchDest_1),
	.datab(temp_branchDest_3),
	.datac(temp_branchDest_2),
	.datad(\Decoder0~30_combout ),
	.cin(gnd),
	.combout(\Decoder0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~32 .lut_mask = 16'h2000;
defparam \Decoder0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N29
dffeas \storeregister[7][1] (
	.clk(!CLK),
	.d(\storeregister[7][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][1] .is_wysiwyg = "true";
defparam \storeregister[7][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N24
cycloneive_lcell_comb \storeregister[6][1]~feeder (
// Equation(s):
// \storeregister[6][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux30),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[6][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[6][1]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[6][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N20
cycloneive_lcell_comb \Decoder0~28 (
// Equation(s):
// \Decoder0~28_combout  = (!temp_branchDest_01 & (temp_regwrite2 & (temp_branchDest_11 & !temp_branchDest_41)))

	.dataa(temp_branchDest_0),
	.datab(temp_regwrite),
	.datac(temp_branchDest_1),
	.datad(temp_branchDest_4),
	.cin(gnd),
	.combout(\Decoder0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~28 .lut_mask = 16'h0040;
defparam \Decoder0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N0
cycloneive_lcell_comb \Decoder0~29 (
// Equation(s):
// \Decoder0~29_combout  = (!temp_branchDest_31 & (\Decoder0~28_combout  & temp_branchDest_21))

	.dataa(temp_branchDest_3),
	.datab(\Decoder0~28_combout ),
	.datac(gnd),
	.datad(temp_branchDest_2),
	.cin(gnd),
	.combout(\Decoder0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~29 .lut_mask = 16'h4400;
defparam \Decoder0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N25
dffeas \storeregister[6][1] (
	.clk(!CLK),
	.d(\storeregister[6][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][1] .is_wysiwyg = "true";
defparam \storeregister[6][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N14
cycloneive_lcell_comb \Mux62~11 (
// Equation(s):
// \Mux62~11_combout  = (\Mux62~10_combout  & (((\storeregister[7][1]~q )) # (!temp_imemload_output_17))) # (!\Mux62~10_combout  & (temp_imemload_output_17 & ((\storeregister[6][1]~q ))))

	.dataa(\Mux62~10_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[7][1]~q ),
	.datad(\storeregister[6][1]~q ),
	.cin(gnd),
	.combout(\Mux62~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~11 .lut_mask = 16'hE6A2;
defparam \Mux62~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N10
cycloneive_lcell_comb \Decoder0~42 (
// Equation(s):
// \Decoder0~42_combout  = (temp_branchDest_11 & (temp_branchDest_31 & (temp_branchDest_21 & \Decoder0~30_combout )))

	.dataa(temp_branchDest_1),
	.datab(temp_branchDest_3),
	.datac(temp_branchDest_2),
	.datad(\Decoder0~30_combout ),
	.cin(gnd),
	.combout(\Decoder0~42_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~42 .lut_mask = 16'h8000;
defparam \Decoder0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y44_N5
dffeas \storeregister[15][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][1] .is_wysiwyg = "true";
defparam \storeregister[15][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N22
cycloneive_lcell_comb \Decoder0~39 (
// Equation(s):
// \Decoder0~39_combout  = (temp_branchDest_21 & (temp_branchDest_31 & \Decoder0~28_combout ))

	.dataa(temp_branchDest_2),
	.datab(temp_branchDest_3),
	.datac(\Decoder0~28_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder0~39_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~39 .lut_mask = 16'h8080;
defparam \Decoder0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N21
dffeas \storeregister[14][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][1] .is_wysiwyg = "true";
defparam \storeregister[14][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N16
cycloneive_lcell_comb \Decoder0~40 (
// Equation(s):
// \Decoder0~40_combout  = (!temp_branchDest_11 & (temp_branchDest_31 & (temp_branchDest_21 & \Decoder0~30_combout )))

	.dataa(temp_branchDest_1),
	.datab(temp_branchDest_3),
	.datac(temp_branchDest_2),
	.datad(\Decoder0~30_combout ),
	.cin(gnd),
	.combout(\Decoder0~40_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~40 .lut_mask = 16'h4000;
defparam \Decoder0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N19
dffeas \storeregister[13][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][1] .is_wysiwyg = "true";
defparam \storeregister[13][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N6
cycloneive_lcell_comb \Decoder0~41 (
// Equation(s):
// \Decoder0~41_combout  = (\Decoder0~18_combout  & (temp_branchDest_21 & !temp_branchDest_41))

	.dataa(\Decoder0~18_combout ),
	.datab(temp_branchDest_2),
	.datac(gnd),
	.datad(temp_branchDest_4),
	.cin(gnd),
	.combout(\Decoder0~41_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~41 .lut_mask = 16'h0088;
defparam \Decoder0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N17
dffeas \storeregister[12][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][1] .is_wysiwyg = "true";
defparam \storeregister[12][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N18
cycloneive_lcell_comb \Mux62~17 (
// Equation(s):
// \Mux62~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[13][1]~q )) # (!temp_imemload_output_16 & ((\storeregister[12][1]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[13][1]~q ),
	.datad(\storeregister[12][1]~q ),
	.cin(gnd),
	.combout(\Mux62~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~17 .lut_mask = 16'hD9C8;
defparam \Mux62~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N26
cycloneive_lcell_comb \Mux62~18 (
// Equation(s):
// \Mux62~18_combout  = (\Mux62~17_combout  & ((\storeregister[15][1]~q ) # ((!temp_imemload_output_17)))) # (!\Mux62~17_combout  & (((\storeregister[14][1]~q  & temp_imemload_output_17))))

	.dataa(\storeregister[15][1]~q ),
	.datab(\storeregister[14][1]~q ),
	.datac(\Mux62~17_combout ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux62~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~18 .lut_mask = 16'hACF0;
defparam \Mux62~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N22
cycloneive_lcell_comb \storeregister[2][1]~feeder (
// Equation(s):
// \storeregister[2][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux30),
	.cin(gnd),
	.combout(\storeregister[2][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[2][1]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[2][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N14
cycloneive_lcell_comb \Decoder0~38 (
// Equation(s):
// \Decoder0~38_combout  = (!temp_branchDest_21 & (!temp_branchDest_31 & \Decoder0~28_combout ))

	.dataa(temp_branchDest_2),
	.datab(temp_branchDest_3),
	.datac(gnd),
	.datad(\Decoder0~28_combout ),
	.cin(gnd),
	.combout(\Decoder0~38_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~38 .lut_mask = 16'h1100;
defparam \Decoder0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N23
dffeas \storeregister[2][1] (
	.clk(!CLK),
	.d(\storeregister[2][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][1] .is_wysiwyg = "true";
defparam \storeregister[2][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N2
cycloneive_lcell_comb \Decoder0~46 (
// Equation(s):
// \Decoder0~46_combout  = (!temp_branchDest_11 & (!temp_branchDest_31 & (!temp_branchDest_21 & \Decoder0~30_combout )))

	.dataa(temp_branchDest_1),
	.datab(temp_branchDest_3),
	.datac(temp_branchDest_2),
	.datad(\Decoder0~30_combout ),
	.cin(gnd),
	.combout(\Decoder0~46_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~46 .lut_mask = 16'h0100;
defparam \Decoder0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N23
dffeas \storeregister[1][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][1] .is_wysiwyg = "true";
defparam \storeregister[1][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N26
cycloneive_lcell_comb \Decoder0~37 (
// Equation(s):
// \Decoder0~37_combout  = (temp_branchDest_11 & (!temp_branchDest_31 & (!temp_branchDest_21 & \Decoder0~30_combout )))

	.dataa(temp_branchDest_1),
	.datab(temp_branchDest_3),
	.datac(temp_branchDest_2),
	.datad(\Decoder0~30_combout ),
	.cin(gnd),
	.combout(\Decoder0~37_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~37 .lut_mask = 16'h0200;
defparam \Decoder0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N13
dffeas \storeregister[3][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][1] .is_wysiwyg = "true";
defparam \storeregister[3][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N22
cycloneive_lcell_comb \Mux62~14 (
// Equation(s):
// \Mux62~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[3][1]~q ))) # (!temp_imemload_output_17 & (\storeregister[1][1]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[1][1]~q ),
	.datad(\storeregister[3][1]~q ),
	.cin(gnd),
	.combout(\Mux62~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~14 .lut_mask = 16'hA820;
defparam \Mux62~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N0
cycloneive_lcell_comb \Mux62~15 (
// Equation(s):
// \Mux62~15_combout  = (\Mux62~14_combout ) # ((!temp_imemload_output_16 & (\storeregister[2][1]~q  & temp_imemload_output_17)))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[2][1]~q ),
	.datac(temp_imemload_output_17),
	.datad(\Mux62~14_combout ),
	.cin(gnd),
	.combout(\Mux62~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~15 .lut_mask = 16'hFF40;
defparam \Mux62~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N16
cycloneive_lcell_comb \storeregister[11][1]~feeder (
// Equation(s):
// \storeregister[11][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux30),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[11][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[11][1]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[11][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N4
cycloneive_lcell_comb \Decoder0~36 (
// Equation(s):
// \Decoder0~36_combout  = (temp_branchDest_11 & (temp_branchDest_31 & (!temp_branchDest_21 & \Decoder0~30_combout )))

	.dataa(temp_branchDest_1),
	.datab(temp_branchDest_3),
	.datac(temp_branchDest_2),
	.datad(\Decoder0~30_combout ),
	.cin(gnd),
	.combout(\Decoder0~36_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~36 .lut_mask = 16'h0800;
defparam \Decoder0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N17
dffeas \storeregister[11][1] (
	.clk(!CLK),
	.d(\storeregister[11][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][1] .is_wysiwyg = "true";
defparam \storeregister[11][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N20
cycloneive_lcell_comb \Decoder0~33 (
// Equation(s):
// \Decoder0~33_combout  = (!temp_branchDest_11 & (temp_branchDest_31 & (!temp_branchDest_21 & \Decoder0~30_combout )))

	.dataa(temp_branchDest_1),
	.datab(temp_branchDest_3),
	.datac(temp_branchDest_2),
	.datad(\Decoder0~30_combout ),
	.cin(gnd),
	.combout(\Decoder0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~33 .lut_mask = 16'h0400;
defparam \Decoder0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N15
dffeas \storeregister[9][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][1] .is_wysiwyg = "true";
defparam \storeregister[9][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N4
cycloneive_lcell_comb \Mux62~13 (
// Equation(s):
// \Mux62~13_combout  = (\Mux62~12_combout  & ((\storeregister[11][1]~q ) # ((!temp_imemload_output_16)))) # (!\Mux62~12_combout  & (((temp_imemload_output_16 & \storeregister[9][1]~q ))))

	.dataa(\Mux62~12_combout ),
	.datab(\storeregister[11][1]~q ),
	.datac(temp_imemload_output_16),
	.datad(\storeregister[9][1]~q ),
	.cin(gnd),
	.combout(\Mux62~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~13 .lut_mask = 16'hDA8A;
defparam \Mux62~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N6
cycloneive_lcell_comb \Mux62~16 (
// Equation(s):
// \Mux62~16_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\Mux62~13_combout ))) # (!temp_imemload_output_19 & (\Mux62~15_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\Mux62~15_combout ),
	.datac(\Mux62~13_combout ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux62~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~16 .lut_mask = 16'hFA44;
defparam \Mux62~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N30
cycloneive_lcell_comb \storeregister[28][1]~feeder (
// Equation(s):
// \storeregister[28][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux30),
	.cin(gnd),
	.combout(\storeregister[28][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][1]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[28][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N30
cycloneive_lcell_comb \Decoder0~23 (
// Equation(s):
// \Decoder0~23_combout  = (\Decoder0~18_combout  & (temp_branchDest_21 & temp_branchDest_41))

	.dataa(\Decoder0~18_combout ),
	.datab(temp_branchDest_2),
	.datac(gnd),
	.datad(temp_branchDest_4),
	.cin(gnd),
	.combout(\Decoder0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~23 .lut_mask = 16'h8800;
defparam \Decoder0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N31
dffeas \storeregister[28][1] (
	.clk(!CLK),
	.d(\storeregister[28][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][1] .is_wysiwyg = "true";
defparam \storeregister[28][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N14
cycloneive_lcell_comb \Mux30~5 (
// Equation(s):
// \Mux30~5_combout  = (\Mux30~4_combout  & (((\storeregister[28][1]~q ) # (!temp_imemload_output_24)))) # (!\Mux30~4_combout  & (\storeregister[24][1]~q  & ((temp_imemload_output_24))))

	.dataa(\Mux30~4_combout ),
	.datab(\storeregister[24][1]~q ),
	.datac(\storeregister[28][1]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~5 .lut_mask = 16'hE4AA;
defparam \Mux30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N14
cycloneive_lcell_comb \Mux30~3 (
// Equation(s):
// \Mux30~3_combout  = (\Mux30~2_combout  & (((\storeregister[30][1]~q )) # (!temp_imemload_output_24))) # (!\Mux30~2_combout  & (temp_imemload_output_24 & (\storeregister[26][1]~q )))

	.dataa(\Mux30~2_combout ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[26][1]~q ),
	.datad(\storeregister[30][1]~q ),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~3 .lut_mask = 16'hEA62;
defparam \Mux30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N12
cycloneive_lcell_comb \Mux30~6 (
// Equation(s):
// \Mux30~6_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & ((\Mux30~3_combout ))) # (!temp_imemload_output_22 & (\Mux30~5_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\Mux30~5_combout ),
	.datad(\Mux30~3_combout ),
	.cin(gnd),
	.combout(\Mux30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~6 .lut_mask = 16'hDC98;
defparam \Mux30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N24
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (temp_imemload_output_24 & ((\storeregister[25][1]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[17][1]~q  & !temp_imemload_output_23))))

	.dataa(\storeregister[25][1]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[17][1]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hCCB8;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N22
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (temp_imemload_output_23 & ((\Mux30~0_combout  & ((\storeregister[29][1]~q ))) # (!\Mux30~0_combout  & (\storeregister[21][1]~q )))) # (!temp_imemload_output_23 & (\Mux30~0_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux30~0_combout ),
	.datac(\storeregister[21][1]~q ),
	.datad(\storeregister[29][1]~q ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hEC64;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N8
cycloneive_lcell_comb \Mux30~7 (
// Equation(s):
// \Mux30~7_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[27][1]~q )) # (!temp_imemload_output_24 & ((\storeregister[19][1]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[27][1]~q ),
	.datad(\storeregister[19][1]~q ),
	.cin(gnd),
	.combout(\Mux30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~7 .lut_mask = 16'hD9C8;
defparam \Mux30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N26
cycloneive_lcell_comb \Mux30~8 (
// Equation(s):
// \Mux30~8_combout  = (\Mux30~7_combout  & ((\storeregister[31][1]~q ) # ((!temp_imemload_output_23)))) # (!\Mux30~7_combout  & (((temp_imemload_output_23 & \storeregister[23][1]~q ))))

	.dataa(\storeregister[31][1]~q ),
	.datab(\Mux30~7_combout ),
	.datac(temp_imemload_output_23),
	.datad(\storeregister[23][1]~q ),
	.cin(gnd),
	.combout(\Mux30~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~8 .lut_mask = 16'hBC8C;
defparam \Mux30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N8
cycloneive_lcell_comb \Decoder0~31 (
// Equation(s):
// \Decoder0~31_combout  = (\Decoder0~20_combout  & (!temp_branchDest_41 & (\Decoder0~8_combout  & temp_branchDest_21)))

	.dataa(\Decoder0~20_combout ),
	.datab(temp_branchDest_4),
	.datac(\Decoder0~8_combout ),
	.datad(temp_branchDest_2),
	.cin(gnd),
	.combout(\Decoder0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~31 .lut_mask = 16'h2000;
defparam \Decoder0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y42_N23
dffeas \storeregister[4][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][1] .is_wysiwyg = "true";
defparam \storeregister[4][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N22
cycloneive_lcell_comb \Mux30~10 (
// Equation(s):
// \Mux30~10_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & (\storeregister[5][1]~q )) # (!temp_imemload_output_21 & ((\storeregister[4][1]~q )))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[5][1]~q ),
	.datac(\storeregister[4][1]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux30~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~10 .lut_mask = 16'hEE50;
defparam \Mux30~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N6
cycloneive_lcell_comb \Mux30~11 (
// Equation(s):
// \Mux30~11_combout  = (\Mux30~10_combout  & (((\storeregister[7][1]~q )) # (!temp_imemload_output_22))) # (!\Mux30~10_combout  & (temp_imemload_output_22 & (\storeregister[6][1]~q )))

	.dataa(\Mux30~10_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[6][1]~q ),
	.datad(\storeregister[7][1]~q ),
	.cin(gnd),
	.combout(\Mux30~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~11 .lut_mask = 16'hEA62;
defparam \Mux30~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N22
cycloneive_lcell_comb \Decoder0~34 (
// Equation(s):
// \Decoder0~34_combout  = (temp_branchDest_31 & (\Decoder0~28_combout  & !temp_branchDest_21))

	.dataa(temp_branchDest_3),
	.datab(\Decoder0~28_combout ),
	.datac(gnd),
	.datad(temp_branchDest_2),
	.cin(gnd),
	.combout(\Decoder0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~34 .lut_mask = 16'h0088;
defparam \Decoder0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N29
dffeas \storeregister[10][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][1] .is_wysiwyg = "true";
defparam \storeregister[10][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N8
cycloneive_lcell_comb \storeregister[8][1]~feeder (
// Equation(s):
// \storeregister[8][1]~feeder_combout  = Mux30

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux30),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[8][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[8][1]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[8][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N0
cycloneive_lcell_comb \Decoder0~18 (
// Equation(s):
// \Decoder0~18_combout  = (!temp_branchDest_01 & (temp_branchDest_31 & (!temp_branchDest_11 & temp_regwrite2)))

	.dataa(temp_branchDest_0),
	.datab(temp_branchDest_3),
	.datac(temp_branchDest_1),
	.datad(temp_regwrite),
	.cin(gnd),
	.combout(\Decoder0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~18 .lut_mask = 16'h0400;
defparam \Decoder0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N22
cycloneive_lcell_comb \Decoder0~35 (
// Equation(s):
// \Decoder0~35_combout  = (!temp_branchDest_41 & (!temp_branchDest_21 & \Decoder0~18_combout ))

	.dataa(temp_branchDest_4),
	.datab(gnd),
	.datac(temp_branchDest_2),
	.datad(\Decoder0~18_combout ),
	.cin(gnd),
	.combout(\Decoder0~35_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~35 .lut_mask = 16'h0500;
defparam \Decoder0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N9
dffeas \storeregister[8][1] (
	.clk(!CLK),
	.d(\storeregister[8][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][1] .is_wysiwyg = "true";
defparam \storeregister[8][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N28
cycloneive_lcell_comb \Mux30~12 (
// Equation(s):
// \Mux30~12_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[10][1]~q )) # (!temp_imemload_output_22 & ((\storeregister[8][1]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][1]~q ),
	.datad(\storeregister[8][1]~q ),
	.cin(gnd),
	.combout(\Mux30~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~12 .lut_mask = 16'hD9C8;
defparam \Mux30~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N14
cycloneive_lcell_comb \Mux30~13 (
// Equation(s):
// \Mux30~13_combout  = (temp_imemload_output_21 & ((\Mux30~12_combout  & (\storeregister[11][1]~q )) # (!\Mux30~12_combout  & ((\storeregister[9][1]~q ))))) # (!temp_imemload_output_21 & (((\Mux30~12_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[11][1]~q ),
	.datac(\storeregister[9][1]~q ),
	.datad(\Mux30~12_combout ),
	.cin(gnd),
	.combout(\Mux30~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~13 .lut_mask = 16'hDDA0;
defparam \Mux30~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N6
cycloneive_lcell_comb \Mux30~15 (
// Equation(s):
// \Mux30~15_combout  = (\Mux30~14_combout ) # ((!temp_imemload_output_21 & (\storeregister[2][1]~q  & temp_imemload_output_22)))

	.dataa(\Mux30~14_combout ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[2][1]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux30~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~15 .lut_mask = 16'hBAAA;
defparam \Mux30~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N28
cycloneive_lcell_comb \Mux30~16 (
// Equation(s):
// \Mux30~16_combout  = (temp_imemload_output_24 & ((\Mux30~13_combout ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((!temp_imemload_output_23 & \Mux30~15_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\Mux30~13_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux30~15_combout ),
	.cin(gnd),
	.combout(\Mux30~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~16 .lut_mask = 16'hADA8;
defparam \Mux30~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N16
cycloneive_lcell_comb \Mux30~17 (
// Equation(s):
// \Mux30~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][1]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[12][1]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[12][1]~q ),
	.datad(\storeregister[13][1]~q ),
	.cin(gnd),
	.combout(\Mux30~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~17 .lut_mask = 16'hBA98;
defparam \Mux30~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N20
cycloneive_lcell_comb \Mux30~18 (
// Equation(s):
// \Mux30~18_combout  = (temp_imemload_output_22 & ((\Mux30~17_combout  & (\storeregister[15][1]~q )) # (!\Mux30~17_combout  & ((\storeregister[14][1]~q ))))) # (!temp_imemload_output_22 & (((\Mux30~17_combout ))))

	.dataa(\storeregister[15][1]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[14][1]~q ),
	.datad(\Mux30~17_combout ),
	.cin(gnd),
	.combout(\Mux30~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~18 .lut_mask = 16'hBBC0;
defparam \Mux30~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N6
cycloneive_lcell_comb \storeregister[29][0]~feeder (
// Equation(s):
// \storeregister[29][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux31),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[29][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][0]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[29][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N7
dffeas \storeregister[29][0] (
	.clk(!CLK),
	.d(\storeregister[29][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][0] .is_wysiwyg = "true";
defparam \storeregister[29][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N0
cycloneive_lcell_comb \storeregister[25][0]~feeder (
// Equation(s):
// \storeregister[25][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux31),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[25][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[25][0]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[25][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N1
dffeas \storeregister[25][0] (
	.clk(!CLK),
	.d(\storeregister[25][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][0] .is_wysiwyg = "true";
defparam \storeregister[25][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N17
dffeas \storeregister[21][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][0] .is_wysiwyg = "true";
defparam \storeregister[21][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N3
dffeas \storeregister[17][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][0] .is_wysiwyg = "true";
defparam \storeregister[17][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N16
cycloneive_lcell_comb \Mux63~0 (
// Equation(s):
// \Mux63~0_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[21][0]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[17][0]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[21][0]~q ),
	.datad(\storeregister[17][0]~q ),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~0 .lut_mask = 16'hB9A8;
defparam \Mux63~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N4
cycloneive_lcell_comb \Mux63~1 (
// Equation(s):
// \Mux63~1_combout  = (\Mux63~0_combout  & ((\storeregister[29][0]~q ) # ((!temp_imemload_output_19)))) # (!\Mux63~0_combout  & (((\storeregister[25][0]~q  & temp_imemload_output_19))))

	.dataa(\storeregister[29][0]~q ),
	.datab(\storeregister[25][0]~q ),
	.datac(\Mux63~0_combout ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~1 .lut_mask = 16'hACF0;
defparam \Mux63~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N3
dffeas \storeregister[30][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][0] .is_wysiwyg = "true";
defparam \storeregister[30][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N26
cycloneive_lcell_comb \Decoder0~15 (
// Equation(s):
// \Decoder0~15_combout  = (\Decoder0~13_combout  & (temp_branchDest_41 & (!temp_branchDest_31 & temp_branchDest_21)))

	.dataa(\Decoder0~13_combout ),
	.datab(temp_branchDest_4),
	.datac(temp_branchDest_3),
	.datad(temp_branchDest_2),
	.cin(gnd),
	.combout(\Decoder0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~15 .lut_mask = 16'h0800;
defparam \Decoder0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N25
dffeas \storeregister[22][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][0] .is_wysiwyg = "true";
defparam \storeregister[22][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N24
cycloneive_lcell_comb \Mux63~3 (
// Equation(s):
// \Mux63~3_combout  = (\Mux63~2_combout  & ((\storeregister[30][0]~q ) # ((!temp_imemload_output_18)))) # (!\Mux63~2_combout  & (((\storeregister[22][0]~q  & temp_imemload_output_18))))

	.dataa(\Mux63~2_combout ),
	.datab(\storeregister[30][0]~q ),
	.datac(\storeregister[22][0]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux63~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~3 .lut_mask = 16'hD8AA;
defparam \Mux63~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N17
dffeas \storeregister[20][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][0] .is_wysiwyg = "true";
defparam \storeregister[20][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N27
dffeas \storeregister[28][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][0] .is_wysiwyg = "true";
defparam \storeregister[28][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N16
cycloneive_lcell_comb \Mux63~5 (
// Equation(s):
// \Mux63~5_combout  = (\Mux63~4_combout  & (((\storeregister[28][0]~q )) # (!temp_imemload_output_18))) # (!\Mux63~4_combout  & (temp_imemload_output_18 & (\storeregister[20][0]~q )))

	.dataa(\Mux63~4_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[20][0]~q ),
	.datad(\storeregister[28][0]~q ),
	.cin(gnd),
	.combout(\Mux63~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~5 .lut_mask = 16'hEA62;
defparam \Mux63~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N0
cycloneive_lcell_comb \Mux63~6 (
// Equation(s):
// \Mux63~6_combout  = (temp_imemload_output_17 & ((\Mux63~3_combout ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((!temp_imemload_output_16 & \Mux63~5_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\Mux63~3_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux63~5_combout ),
	.cin(gnd),
	.combout(\Mux63~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~6 .lut_mask = 16'hADA8;
defparam \Mux63~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N22
cycloneive_lcell_comb \storeregister[23][0]~feeder (
// Equation(s):
// \storeregister[23][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux31),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[23][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][0]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[23][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N23
dffeas \storeregister[23][0] (
	.clk(!CLK),
	.d(\storeregister[23][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][0] .is_wysiwyg = "true";
defparam \storeregister[23][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N12
cycloneive_lcell_comb \Mux63~7 (
// Equation(s):
// \Mux63~7_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[23][0]~q ))) # (!temp_imemload_output_18 & (\storeregister[19][0]~q ))))

	.dataa(\storeregister[19][0]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[23][0]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux63~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~7 .lut_mask = 16'hFC22;
defparam \Mux63~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N2
cycloneive_lcell_comb \storeregister[27][0]~feeder (
// Equation(s):
// \storeregister[27][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux31),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][0]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N3
dffeas \storeregister[27][0] (
	.clk(!CLK),
	.d(\storeregister[27][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][0] .is_wysiwyg = "true";
defparam \storeregister[27][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N4
cycloneive_lcell_comb \storeregister[31][0]~feeder (
// Equation(s):
// \storeregister[31][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux31),
	.cin(gnd),
	.combout(\storeregister[31][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][0]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[31][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N5
dffeas \storeregister[31][0] (
	.clk(!CLK),
	.d(\storeregister[31][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][0] .is_wysiwyg = "true";
defparam \storeregister[31][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N14
cycloneive_lcell_comb \Mux63~8 (
// Equation(s):
// \Mux63~8_combout  = (\Mux63~7_combout  & (((\storeregister[31][0]~q ) # (!temp_imemload_output_19)))) # (!\Mux63~7_combout  & (\storeregister[27][0]~q  & ((temp_imemload_output_19))))

	.dataa(\Mux63~7_combout ),
	.datab(\storeregister[27][0]~q ),
	.datac(\storeregister[31][0]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux63~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~8 .lut_mask = 16'hE4AA;
defparam \Mux63~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N13
dffeas \storeregister[10][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][0] .is_wysiwyg = "true";
defparam \storeregister[10][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N24
cycloneive_lcell_comb \Mux63~10 (
// Equation(s):
// \Mux63~10_combout  = (temp_imemload_output_17 & (((\storeregister[10][0]~q ) # (temp_imemload_output_16)))) # (!temp_imemload_output_17 & (\storeregister[8][0]~q  & ((!temp_imemload_output_16))))

	.dataa(\storeregister[8][0]~q ),
	.datab(\storeregister[10][0]~q ),
	.datac(temp_imemload_output_17),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux63~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~10 .lut_mask = 16'hF0CA;
defparam \Mux63~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N3
dffeas \storeregister[11][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][0] .is_wysiwyg = "true";
defparam \storeregister[11][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N7
dffeas \storeregister[9][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][0] .is_wysiwyg = "true";
defparam \storeregister[9][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N2
cycloneive_lcell_comb \Mux63~11 (
// Equation(s):
// \Mux63~11_combout  = (temp_imemload_output_16 & ((\Mux63~10_combout  & (\storeregister[11][0]~q )) # (!\Mux63~10_combout  & ((\storeregister[9][0]~q ))))) # (!temp_imemload_output_16 & (\Mux63~10_combout ))

	.dataa(temp_imemload_output_16),
	.datab(\Mux63~10_combout ),
	.datac(\storeregister[11][0]~q ),
	.datad(\storeregister[9][0]~q ),
	.cin(gnd),
	.combout(\Mux63~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~11 .lut_mask = 16'hE6C4;
defparam \Mux63~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N16
cycloneive_lcell_comb \storeregister[6][0]~feeder (
// Equation(s):
// \storeregister[6][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux31),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[6][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[6][0]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[6][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N17
dffeas \storeregister[6][0] (
	.clk(!CLK),
	.d(\storeregister[6][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][0] .is_wysiwyg = "true";
defparam \storeregister[6][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N0
cycloneive_lcell_comb \storeregister[7][0]~feeder (
// Equation(s):
// \storeregister[7][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux31),
	.cin(gnd),
	.combout(\storeregister[7][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[7][0]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[7][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N1
dffeas \storeregister[7][0] (
	.clk(!CLK),
	.d(\storeregister[7][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][0] .is_wysiwyg = "true";
defparam \storeregister[7][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N22
cycloneive_lcell_comb \Mux63~13 (
// Equation(s):
// \Mux63~13_combout  = (\Mux63~12_combout  & (((\storeregister[7][0]~q ) # (!temp_imemload_output_17)))) # (!\Mux63~12_combout  & (\storeregister[6][0]~q  & (temp_imemload_output_17)))

	.dataa(\Mux63~12_combout ),
	.datab(\storeregister[6][0]~q ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[7][0]~q ),
	.cin(gnd),
	.combout(\Mux63~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~13 .lut_mask = 16'hEA4A;
defparam \Mux63~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N25
dffeas \storeregister[2][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][0] .is_wysiwyg = "true";
defparam \storeregister[2][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N18
cycloneive_lcell_comb \Mux63~15 (
// Equation(s):
// \Mux63~15_combout  = (\Mux63~14_combout ) # ((\storeregister[2][0]~q  & (temp_imemload_output_17 & !temp_imemload_output_16)))

	.dataa(\Mux63~14_combout ),
	.datab(\storeregister[2][0]~q ),
	.datac(temp_imemload_output_17),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux63~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~15 .lut_mask = 16'hAAEA;
defparam \Mux63~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N4
cycloneive_lcell_comb \Mux63~16 (
// Equation(s):
// \Mux63~16_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\Mux63~13_combout )) # (!temp_imemload_output_18 & ((\Mux63~15_combout )))))

	.dataa(temp_imemload_output_19),
	.datab(\Mux63~13_combout ),
	.datac(\Mux63~15_combout ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux63~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~16 .lut_mask = 16'hEE50;
defparam \Mux63~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N4
cycloneive_lcell_comb \storeregister[15][0]~feeder (
// Equation(s):
// \storeregister[15][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux31),
	.cin(gnd),
	.combout(\storeregister[15][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][0]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y44_N5
dffeas \storeregister[15][0] (
	.clk(!CLK),
	.d(\storeregister[15][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][0] .is_wysiwyg = "true";
defparam \storeregister[15][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N20
cycloneive_lcell_comb \storeregister[12][0]~feeder (
// Equation(s):
// \storeregister[12][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux31),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[12][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[12][0]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[12][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N21
dffeas \storeregister[12][0] (
	.clk(!CLK),
	.d(\storeregister[12][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][0] .is_wysiwyg = "true";
defparam \storeregister[12][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N0
cycloneive_lcell_comb \storeregister[13][0]~feeder (
// Equation(s):
// \storeregister[13][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux31),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[13][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[13][0]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[13][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N1
dffeas \storeregister[13][0] (
	.clk(!CLK),
	.d(\storeregister[13][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][0] .is_wysiwyg = "true";
defparam \storeregister[13][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N18
cycloneive_lcell_comb \Mux63~17 (
// Equation(s):
// \Mux63~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][0]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][0]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[12][0]~q ),
	.datad(\storeregister[13][0]~q ),
	.cin(gnd),
	.combout(\Mux63~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~17 .lut_mask = 16'hDC98;
defparam \Mux63~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N2
cycloneive_lcell_comb \storeregister[14][0]~feeder (
// Equation(s):
// \storeregister[14][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux31),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[14][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][0]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[14][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N3
dffeas \storeregister[14][0] (
	.clk(!CLK),
	.d(\storeregister[14][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][0] .is_wysiwyg = "true";
defparam \storeregister[14][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N8
cycloneive_lcell_comb \Mux63~18 (
// Equation(s):
// \Mux63~18_combout  = (temp_imemload_output_17 & ((\Mux63~17_combout  & (\storeregister[15][0]~q )) # (!\Mux63~17_combout  & ((\storeregister[14][0]~q ))))) # (!temp_imemload_output_17 & (((\Mux63~17_combout ))))

	.dataa(\storeregister[15][0]~q ),
	.datab(temp_imemload_output_17),
	.datac(\Mux63~17_combout ),
	.datad(\storeregister[14][0]~q ),
	.cin(gnd),
	.combout(\Mux63~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~18 .lut_mask = 16'hBCB0;
defparam \Mux63~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N2
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[21][0]~q )) # (!temp_imemload_output_23 & ((\storeregister[17][0]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[21][0]~q ),
	.datac(\storeregister[17][0]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'hEE50;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N12
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (temp_imemload_output_24 & ((\Mux31~0_combout  & (\storeregister[29][0]~q )) # (!\Mux31~0_combout  & ((\storeregister[25][0]~q ))))) # (!temp_imemload_output_24 & (\Mux31~0_combout ))

	.dataa(temp_imemload_output_24),
	.datab(\Mux31~0_combout ),
	.datac(\storeregister[29][0]~q ),
	.datad(\storeregister[25][0]~q ),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hE6C4;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N30
cycloneive_lcell_comb \storeregister[19][0]~feeder (
// Equation(s):
// \storeregister[19][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux31),
	.cin(gnd),
	.combout(\storeregister[19][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[19][0]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[19][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N31
dffeas \storeregister[19][0] (
	.clk(!CLK),
	.d(\storeregister[19][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][0] .is_wysiwyg = "true";
defparam \storeregister[19][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N14
cycloneive_lcell_comb \Mux31~7 (
// Equation(s):
// \Mux31~7_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[23][0]~q ))) # (!temp_imemload_output_23 & (\storeregister[19][0]~q ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[19][0]~q ),
	.datac(\storeregister[23][0]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~7 .lut_mask = 16'hFA44;
defparam \Mux31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N28
cycloneive_lcell_comb \Mux31~8 (
// Equation(s):
// \Mux31~8_combout  = (temp_imemload_output_24 & ((\Mux31~7_combout  & (\storeregister[31][0]~q )) # (!\Mux31~7_combout  & ((\storeregister[27][0]~q ))))) # (!temp_imemload_output_24 & (((\Mux31~7_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[31][0]~q ),
	.datac(\Mux31~7_combout ),
	.datad(\storeregister[27][0]~q ),
	.cin(gnd),
	.combout(\Mux31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~8 .lut_mask = 16'hDAD0;
defparam \Mux31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N29
dffeas \storeregister[24][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][0] .is_wysiwyg = "true";
defparam \storeregister[24][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N31
dffeas \storeregister[16][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][0] .is_wysiwyg = "true";
defparam \storeregister[16][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N28
cycloneive_lcell_comb \Mux31~4 (
// Equation(s):
// \Mux31~4_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[24][0]~q )) # (!temp_imemload_output_24 & ((\storeregister[16][0]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[24][0]~q ),
	.datad(\storeregister[16][0]~q ),
	.cin(gnd),
	.combout(\Mux31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~4 .lut_mask = 16'hD9C8;
defparam \Mux31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N26
cycloneive_lcell_comb \Mux31~5 (
// Equation(s):
// \Mux31~5_combout  = (temp_imemload_output_23 & ((\Mux31~4_combout  & ((\storeregister[28][0]~q ))) # (!\Mux31~4_combout  & (\storeregister[20][0]~q )))) # (!temp_imemload_output_23 & (((\Mux31~4_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[20][0]~q ),
	.datac(\storeregister[28][0]~q ),
	.datad(\Mux31~4_combout ),
	.cin(gnd),
	.combout(\Mux31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~5 .lut_mask = 16'hF588;
defparam \Mux31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N2
cycloneive_lcell_comb \Mux31~3 (
// Equation(s):
// \Mux31~3_combout  = (\Mux31~2_combout  & (((\storeregister[30][0]~q )) # (!temp_imemload_output_23))) # (!\Mux31~2_combout  & (temp_imemload_output_23 & ((\storeregister[22][0]~q ))))

	.dataa(\Mux31~2_combout ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[30][0]~q ),
	.datad(\storeregister[22][0]~q ),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~3 .lut_mask = 16'hE6A2;
defparam \Mux31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N4
cycloneive_lcell_comb \Mux31~6 (
// Equation(s):
// \Mux31~6_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21) # (\Mux31~3_combout )))) # (!temp_imemload_output_22 & (\Mux31~5_combout  & (!temp_imemload_output_21)))

	.dataa(\Mux31~5_combout ),
	.datab(temp_imemload_output_22),
	.datac(temp_imemload_output_21),
	.datad(\Mux31~3_combout ),
	.cin(gnd),
	.combout(\Mux31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~6 .lut_mask = 16'hCEC2;
defparam \Mux31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N17
dffeas \storeregister[3][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][0] .is_wysiwyg = "true";
defparam \storeregister[3][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N16
cycloneive_lcell_comb \Mux31~14 (
// Equation(s):
// \Mux31~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][0]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][0]~q ))))

	.dataa(\storeregister[1][0]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[3][0]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux31~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~14 .lut_mask = 16'hE200;
defparam \Mux31~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N24
cycloneive_lcell_comb \Mux31~15 (
// Equation(s):
// \Mux31~15_combout  = (\Mux31~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][0]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][0]~q ),
	.datad(\Mux31~14_combout ),
	.cin(gnd),
	.combout(\Mux31~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~15 .lut_mask = 16'hFF40;
defparam \Mux31~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y42_N17
dffeas \storeregister[5][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][0] .is_wysiwyg = "true";
defparam \storeregister[5][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y42_N15
dffeas \storeregister[4][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][0] .is_wysiwyg = "true";
defparam \storeregister[4][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N14
cycloneive_lcell_comb \Mux31~12 (
// Equation(s):
// \Mux31~12_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & (\storeregister[5][0]~q )) # (!temp_imemload_output_21 & ((\storeregister[4][0]~q )))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[5][0]~q ),
	.datac(\storeregister[4][0]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux31~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~12 .lut_mask = 16'hEE50;
defparam \Mux31~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N20
cycloneive_lcell_comb \Mux31~13 (
// Equation(s):
// \Mux31~13_combout  = (temp_imemload_output_22 & ((\Mux31~12_combout  & (\storeregister[7][0]~q )) # (!\Mux31~12_combout  & ((\storeregister[6][0]~q ))))) # (!temp_imemload_output_22 & (((\Mux31~12_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[7][0]~q ),
	.datac(\Mux31~12_combout ),
	.datad(\storeregister[6][0]~q ),
	.cin(gnd),
	.combout(\Mux31~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~13 .lut_mask = 16'hDAD0;
defparam \Mux31~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N10
cycloneive_lcell_comb \Mux31~16 (
// Equation(s):
// \Mux31~16_combout  = (temp_imemload_output_23 & (((\Mux31~13_combout ) # (temp_imemload_output_24)))) # (!temp_imemload_output_23 & (\Mux31~15_combout  & ((!temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\Mux31~15_combout ),
	.datac(\Mux31~13_combout ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux31~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~16 .lut_mask = 16'hAAE4;
defparam \Mux31~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N10
cycloneive_lcell_comb \storeregister[8][0]~feeder (
// Equation(s):
// \storeregister[8][0]~feeder_combout  = Mux31

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux31),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[8][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[8][0]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[8][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N11
dffeas \storeregister[8][0] (
	.clk(!CLK),
	.d(\storeregister[8][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][0] .is_wysiwyg = "true";
defparam \storeregister[8][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N12
cycloneive_lcell_comb \Mux31~10 (
// Equation(s):
// \Mux31~10_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[10][0]~q )) # (!temp_imemload_output_22 & ((\storeregister[8][0]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][0]~q ),
	.datad(\storeregister[8][0]~q ),
	.cin(gnd),
	.combout(\Mux31~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~10 .lut_mask = 16'hD9C8;
defparam \Mux31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N6
cycloneive_lcell_comb \Mux31~11 (
// Equation(s):
// \Mux31~11_combout  = (temp_imemload_output_21 & ((\Mux31~10_combout  & ((\storeregister[11][0]~q ))) # (!\Mux31~10_combout  & (\storeregister[9][0]~q )))) # (!temp_imemload_output_21 & (\Mux31~10_combout ))

	.dataa(temp_imemload_output_21),
	.datab(\Mux31~10_combout ),
	.datac(\storeregister[9][0]~q ),
	.datad(\storeregister[11][0]~q ),
	.cin(gnd),
	.combout(\Mux31~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~11 .lut_mask = 16'hEC64;
defparam \Mux31~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N24
cycloneive_lcell_comb \Mux31~17 (
// Equation(s):
// \Mux31~17_combout  = (temp_imemload_output_21 & ((\storeregister[13][0]~q ) # ((temp_imemload_output_22)))) # (!temp_imemload_output_21 & (((\storeregister[12][0]~q  & !temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[13][0]~q ),
	.datac(\storeregister[12][0]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux31~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~17 .lut_mask = 16'hAAD8;
defparam \Mux31~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N8
cycloneive_lcell_comb \Mux31~18 (
// Equation(s):
// \Mux31~18_combout  = (\Mux31~17_combout  & (((\storeregister[15][0]~q ) # (!temp_imemload_output_22)))) # (!\Mux31~17_combout  & (\storeregister[14][0]~q  & (temp_imemload_output_22)))

	.dataa(\storeregister[14][0]~q ),
	.datab(\Mux31~17_combout ),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[15][0]~q ),
	.cin(gnd),
	.combout(\Mux31~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~18 .lut_mask = 16'hEC2C;
defparam \Mux31~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N1
dffeas \storeregister[20][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][2] .is_wysiwyg = "true";
defparam \storeregister[20][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N23
dffeas \storeregister[16][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][2] .is_wysiwyg = "true";
defparam \storeregister[16][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N8
cycloneive_lcell_comb \storeregister[24][2]~feeder (
// Equation(s):
// \storeregister[24][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux29),
	.cin(gnd),
	.combout(\storeregister[24][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][2]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[24][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N9
dffeas \storeregister[24][2] (
	.clk(!CLK),
	.d(\storeregister[24][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][2] .is_wysiwyg = "true";
defparam \storeregister[24][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N22
cycloneive_lcell_comb \Mux29~4 (
// Equation(s):
// \Mux29~4_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[24][2]~q ))) # (!temp_imemload_output_24 & (\storeregister[16][2]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][2]~q ),
	.datad(\storeregister[24][2]~q ),
	.cin(gnd),
	.combout(\Mux29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~4 .lut_mask = 16'hDC98;
defparam \Mux29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N8
cycloneive_lcell_comb \Mux29~5 (
// Equation(s):
// \Mux29~5_combout  = (\Mux29~4_combout  & ((\storeregister[28][2]~q ) # ((!temp_imemload_output_23)))) # (!\Mux29~4_combout  & (((\storeregister[20][2]~q  & temp_imemload_output_23))))

	.dataa(\storeregister[28][2]~q ),
	.datab(\storeregister[20][2]~q ),
	.datac(\Mux29~4_combout ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~5 .lut_mask = 16'hACF0;
defparam \Mux29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N24
cycloneive_lcell_comb \storeregister[30][2]~feeder (
// Equation(s):
// \storeregister[30][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux29),
	.cin(gnd),
	.combout(\storeregister[30][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][2]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[30][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N25
dffeas \storeregister[30][2] (
	.clk(!CLK),
	.d(\storeregister[30][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][2] .is_wysiwyg = "true";
defparam \storeregister[30][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N24
cycloneive_lcell_comb \storeregister[18][2]~feeder (
// Equation(s):
// \storeregister[18][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux29),
	.cin(gnd),
	.combout(\storeregister[18][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[18][2]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[18][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N0
cycloneive_lcell_comb \Decoder0~16 (
// Equation(s):
// \Decoder0~16_combout  = (\Decoder0~13_combout  & (temp_branchDest_41 & (!temp_branchDest_31 & !temp_branchDest_21)))

	.dataa(\Decoder0~13_combout ),
	.datab(temp_branchDest_4),
	.datac(temp_branchDest_3),
	.datad(temp_branchDest_2),
	.cin(gnd),
	.combout(\Decoder0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~16 .lut_mask = 16'h0008;
defparam \Decoder0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N25
dffeas \storeregister[18][2] (
	.clk(!CLK),
	.d(\storeregister[18][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][2] .is_wysiwyg = "true";
defparam \storeregister[18][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N9
dffeas \storeregister[26][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][2] .is_wysiwyg = "true";
defparam \storeregister[26][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N8
cycloneive_lcell_comb \Mux29~2 (
// Equation(s):
// \Mux29~2_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[26][2]~q ))) # (!temp_imemload_output_24 & (\storeregister[18][2]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[18][2]~q ),
	.datac(\storeregister[26][2]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~2 .lut_mask = 16'hFA44;
defparam \Mux29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N2
cycloneive_lcell_comb \Mux29~3 (
// Equation(s):
// \Mux29~3_combout  = (temp_imemload_output_23 & ((\Mux29~2_combout  & ((\storeregister[30][2]~q ))) # (!\Mux29~2_combout  & (\storeregister[22][2]~q )))) # (!temp_imemload_output_23 & (((\Mux29~2_combout ))))

	.dataa(\storeregister[22][2]~q ),
	.datab(\storeregister[30][2]~q ),
	.datac(temp_imemload_output_23),
	.datad(\Mux29~2_combout ),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~3 .lut_mask = 16'hCFA0;
defparam \Mux29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N26
cycloneive_lcell_comb \Mux29~6 (
// Equation(s):
// \Mux29~6_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21) # (\Mux29~3_combout )))) # (!temp_imemload_output_22 & (\Mux29~5_combout  & (!temp_imemload_output_21)))

	.dataa(temp_imemload_output_22),
	.datab(\Mux29~5_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux29~3_combout ),
	.cin(gnd),
	.combout(\Mux29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~6 .lut_mask = 16'hAEA4;
defparam \Mux29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N5
dffeas \storeregister[19][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][2] .is_wysiwyg = "true";
defparam \storeregister[19][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N27
dffeas \storeregister[23][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][2] .is_wysiwyg = "true";
defparam \storeregister[23][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N26
cycloneive_lcell_comb \Mux29~7 (
// Equation(s):
// \Mux29~7_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[23][2]~q ))) # (!temp_imemload_output_23 & (\storeregister[19][2]~q ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[19][2]~q ),
	.datac(\storeregister[23][2]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~7 .lut_mask = 16'hFA44;
defparam \Mux29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N14
cycloneive_lcell_comb \storeregister[31][2]~feeder (
// Equation(s):
// \storeregister[31][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux29),
	.cin(gnd),
	.combout(\storeregister[31][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][2]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[31][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N15
dffeas \storeregister[31][2] (
	.clk(!CLK),
	.d(\storeregister[31][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][2] .is_wysiwyg = "true";
defparam \storeregister[31][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N10
cycloneive_lcell_comb \storeregister[27][2]~feeder (
// Equation(s):
// \storeregister[27][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux29),
	.cin(gnd),
	.combout(\storeregister[27][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][2]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[27][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N11
dffeas \storeregister[27][2] (
	.clk(!CLK),
	.d(\storeregister[27][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][2] .is_wysiwyg = "true";
defparam \storeregister[27][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N4
cycloneive_lcell_comb \Mux29~8 (
// Equation(s):
// \Mux29~8_combout  = (temp_imemload_output_24 & ((\Mux29~7_combout  & (\storeregister[31][2]~q )) # (!\Mux29~7_combout  & ((\storeregister[27][2]~q ))))) # (!temp_imemload_output_24 & (\Mux29~7_combout ))

	.dataa(temp_imemload_output_24),
	.datab(\Mux29~7_combout ),
	.datac(\storeregister[31][2]~q ),
	.datad(\storeregister[27][2]~q ),
	.cin(gnd),
	.combout(\Mux29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~8 .lut_mask = 16'hE6C4;
defparam \Mux29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N3
dffeas \storeregister[25][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][2] .is_wysiwyg = "true";
defparam \storeregister[25][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N1
dffeas \storeregister[29][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][2] .is_wysiwyg = "true";
defparam \storeregister[29][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N21
dffeas \storeregister[17][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][2] .is_wysiwyg = "true";
defparam \storeregister[17][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N20
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[21][2]~q )) # (!temp_imemload_output_23 & ((\storeregister[17][2]~q )))))

	.dataa(\storeregister[21][2]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[17][2]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hEE30;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N0
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (temp_imemload_output_24 & ((\Mux29~0_combout  & ((\storeregister[29][2]~q ))) # (!\Mux29~0_combout  & (\storeregister[25][2]~q )))) # (!temp_imemload_output_24 & (((\Mux29~0_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[25][2]~q ),
	.datac(\storeregister[29][2]~q ),
	.datad(\Mux29~0_combout ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hF588;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y42_N29
dffeas \storeregister[5][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][2] .is_wysiwyg = "true";
defparam \storeregister[5][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y42_N27
dffeas \storeregister[4][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][2] .is_wysiwyg = "true";
defparam \storeregister[4][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N26
cycloneive_lcell_comb \Mux29~12 (
// Equation(s):
// \Mux29~12_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & (\storeregister[5][2]~q )) # (!temp_imemload_output_21 & ((\storeregister[4][2]~q )))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[5][2]~q ),
	.datac(\storeregister[4][2]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux29~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~12 .lut_mask = 16'hEE50;
defparam \Mux29~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N10
cycloneive_lcell_comb \storeregister[6][2]~feeder (
// Equation(s):
// \storeregister[6][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux29),
	.cin(gnd),
	.combout(\storeregister[6][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[6][2]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[6][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N11
dffeas \storeregister[6][2] (
	.clk(!CLK),
	.d(\storeregister[6][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][2] .is_wysiwyg = "true";
defparam \storeregister[6][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N28
cycloneive_lcell_comb \Mux29~13 (
// Equation(s):
// \Mux29~13_combout  = (\Mux29~12_combout  & ((\storeregister[7][2]~q ) # ((!temp_imemload_output_22)))) # (!\Mux29~12_combout  & (((\storeregister[6][2]~q  & temp_imemload_output_22))))

	.dataa(\storeregister[7][2]~q ),
	.datab(\Mux29~12_combout ),
	.datac(\storeregister[6][2]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux29~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~13 .lut_mask = 16'hB8CC;
defparam \Mux29~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N5
dffeas \storeregister[3][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][2] .is_wysiwyg = "true";
defparam \storeregister[3][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N19
dffeas \storeregister[1][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][2] .is_wysiwyg = "true";
defparam \storeregister[1][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N18
cycloneive_lcell_comb \Mux29~14 (
// Equation(s):
// \Mux29~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[3][2]~q )) # (!temp_imemload_output_22 & ((\storeregister[1][2]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[3][2]~q ),
	.datac(\storeregister[1][2]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux29~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~14 .lut_mask = 16'h88A0;
defparam \Mux29~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N18
cycloneive_lcell_comb \Mux29~15 (
// Equation(s):
// \Mux29~15_combout  = (\Mux29~14_combout ) # ((\storeregister[2][2]~q  & (temp_imemload_output_22 & !temp_imemload_output_21)))

	.dataa(\storeregister[2][2]~q ),
	.datab(\Mux29~14_combout ),
	.datac(temp_imemload_output_22),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux29~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~15 .lut_mask = 16'hCCEC;
defparam \Mux29~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N16
cycloneive_lcell_comb \Mux29~16 (
// Equation(s):
// \Mux29~16_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\Mux29~13_combout )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & ((\Mux29~15_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\Mux29~13_combout ),
	.datad(\Mux29~15_combout ),
	.cin(gnd),
	.combout(\Mux29~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~16 .lut_mask = 16'hB9A8;
defparam \Mux29~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N3
dffeas \storeregister[12][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][2] .is_wysiwyg = "true";
defparam \storeregister[12][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N29
dffeas \storeregister[13][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][2] .is_wysiwyg = "true";
defparam \storeregister[13][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N28
cycloneive_lcell_comb \Mux29~17 (
// Equation(s):
// \Mux29~17_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[13][2]~q ))) # (!temp_imemload_output_21 & (\storeregister[12][2]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[12][2]~q ),
	.datac(\storeregister[13][2]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux29~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~17 .lut_mask = 16'hFA44;
defparam \Mux29~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N24
cycloneive_lcell_comb \storeregister[14][2]~feeder (
// Equation(s):
// \storeregister[14][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux29),
	.cin(gnd),
	.combout(\storeregister[14][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][2]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y39_N25
dffeas \storeregister[14][2] (
	.clk(!CLK),
	.d(\storeregister[14][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][2] .is_wysiwyg = "true";
defparam \storeregister[14][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N0
cycloneive_lcell_comb \storeregister[15][2]~feeder (
// Equation(s):
// \storeregister[15][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux29),
	.cin(gnd),
	.combout(\storeregister[15][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][2]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N1
dffeas \storeregister[15][2] (
	.clk(!CLK),
	.d(\storeregister[15][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][2] .is_wysiwyg = "true";
defparam \storeregister[15][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N2
cycloneive_lcell_comb \Mux29~18 (
// Equation(s):
// \Mux29~18_combout  = (\Mux29~17_combout  & (((\storeregister[15][2]~q ) # (!temp_imemload_output_22)))) # (!\Mux29~17_combout  & (\storeregister[14][2]~q  & (temp_imemload_output_22)))

	.dataa(\Mux29~17_combout ),
	.datab(\storeregister[14][2]~q ),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[15][2]~q ),
	.cin(gnd),
	.combout(\Mux29~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~18 .lut_mask = 16'hEA4A;
defparam \Mux29~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N19
dffeas \storeregister[9][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][2] .is_wysiwyg = "true";
defparam \storeregister[9][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N23
dffeas \storeregister[10][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][2] .is_wysiwyg = "true";
defparam \storeregister[10][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N0
cycloneive_lcell_comb \storeregister[8][2]~feeder (
// Equation(s):
// \storeregister[8][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux29),
	.cin(gnd),
	.combout(\storeregister[8][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[8][2]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[8][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N1
dffeas \storeregister[8][2] (
	.clk(!CLK),
	.d(\storeregister[8][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][2] .is_wysiwyg = "true";
defparam \storeregister[8][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N22
cycloneive_lcell_comb \Mux29~10 (
// Equation(s):
// \Mux29~10_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[10][2]~q )) # (!temp_imemload_output_22 & ((\storeregister[8][2]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][2]~q ),
	.datad(\storeregister[8][2]~q ),
	.cin(gnd),
	.combout(\Mux29~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~10 .lut_mask = 16'hD9C8;
defparam \Mux29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N25
dffeas \storeregister[11][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][2] .is_wysiwyg = "true";
defparam \storeregister[11][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N24
cycloneive_lcell_comb \Mux29~11 (
// Equation(s):
// \Mux29~11_combout  = (\Mux29~10_combout  & (((\storeregister[11][2]~q ) # (!temp_imemload_output_21)))) # (!\Mux29~10_combout  & (\storeregister[9][2]~q  & ((temp_imemload_output_21))))

	.dataa(\storeregister[9][2]~q ),
	.datab(\Mux29~10_combout ),
	.datac(\storeregister[11][2]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux29~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~11 .lut_mask = 16'hE2CC;
defparam \Mux29~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N0
cycloneive_lcell_comb \storeregister[31][4]~feeder (
// Equation(s):
// \storeregister[31][4]~feeder_combout  = Mux27

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux27),
	.cin(gnd),
	.combout(\storeregister[31][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][4]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[31][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N1
dffeas \storeregister[31][4] (
	.clk(!CLK),
	.d(\storeregister[31][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][4] .is_wysiwyg = "true";
defparam \storeregister[31][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N15
dffeas \storeregister[27][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][4] .is_wysiwyg = "true";
defparam \storeregister[27][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N31
dffeas \storeregister[23][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][4] .is_wysiwyg = "true";
defparam \storeregister[23][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N17
dffeas \storeregister[19][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][4] .is_wysiwyg = "true";
defparam \storeregister[19][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N30
cycloneive_lcell_comb \Mux27~7 (
// Equation(s):
// \Mux27~7_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[23][4]~q )) # (!temp_imemload_output_23 & ((\storeregister[19][4]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[23][4]~q ),
	.datad(\storeregister[19][4]~q ),
	.cin(gnd),
	.combout(\Mux27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~7 .lut_mask = 16'hD9C8;
defparam \Mux27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N14
cycloneive_lcell_comb \Mux27~8 (
// Equation(s):
// \Mux27~8_combout  = (temp_imemload_output_24 & ((\Mux27~7_combout  & (\storeregister[31][4]~q )) # (!\Mux27~7_combout  & ((\storeregister[27][4]~q ))))) # (!temp_imemload_output_24 & (((\Mux27~7_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[31][4]~q ),
	.datac(\storeregister[27][4]~q ),
	.datad(\Mux27~7_combout ),
	.cin(gnd),
	.combout(\Mux27~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~8 .lut_mask = 16'hDDA0;
defparam \Mux27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N7
dffeas \storeregister[16][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][4] .is_wysiwyg = "true";
defparam \storeregister[16][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N18
cycloneive_lcell_comb \storeregister[24][4]~feeder (
// Equation(s):
// \storeregister[24][4]~feeder_combout  = Mux27

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux27),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[24][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][4]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[24][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N19
dffeas \storeregister[24][4] (
	.clk(!CLK),
	.d(\storeregister[24][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][4] .is_wysiwyg = "true";
defparam \storeregister[24][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N6
cycloneive_lcell_comb \Mux27~4 (
// Equation(s):
// \Mux27~4_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[24][4]~q ))) # (!temp_imemload_output_24 & (\storeregister[16][4]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][4]~q ),
	.datad(\storeregister[24][4]~q ),
	.cin(gnd),
	.combout(\Mux27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~4 .lut_mask = 16'hDC98;
defparam \Mux27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N13
dffeas \storeregister[20][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][4] .is_wysiwyg = "true";
defparam \storeregister[20][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N1
dffeas \storeregister[28][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][4] .is_wysiwyg = "true";
defparam \storeregister[28][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N18
cycloneive_lcell_comb \Mux27~5 (
// Equation(s):
// \Mux27~5_combout  = (temp_imemload_output_23 & ((\Mux27~4_combout  & ((\storeregister[28][4]~q ))) # (!\Mux27~4_combout  & (\storeregister[20][4]~q )))) # (!temp_imemload_output_23 & (\Mux27~4_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux27~4_combout ),
	.datac(\storeregister[20][4]~q ),
	.datad(\storeregister[28][4]~q ),
	.cin(gnd),
	.combout(\Mux27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~5 .lut_mask = 16'hEC64;
defparam \Mux27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N17
dffeas \storeregister[26][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][4] .is_wysiwyg = "true";
defparam \storeregister[26][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N22
cycloneive_lcell_comb \storeregister[18][4]~feeder (
// Equation(s):
// \storeregister[18][4]~feeder_combout  = Mux27

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux27),
	.cin(gnd),
	.combout(\storeregister[18][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[18][4]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[18][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N23
dffeas \storeregister[18][4] (
	.clk(!CLK),
	.d(\storeregister[18][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][4] .is_wysiwyg = "true";
defparam \storeregister[18][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N16
cycloneive_lcell_comb \Mux27~2 (
// Equation(s):
// \Mux27~2_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[26][4]~q )) # (!temp_imemload_output_24 & ((\storeregister[18][4]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[26][4]~q ),
	.datad(\storeregister[18][4]~q ),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~2 .lut_mask = 16'hD9C8;
defparam \Mux27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N11
dffeas \storeregister[22][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][4] .is_wysiwyg = "true";
defparam \storeregister[22][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N6
cycloneive_lcell_comb \storeregister[30][4]~feeder (
// Equation(s):
// \storeregister[30][4]~feeder_combout  = Mux27

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux27),
	.cin(gnd),
	.combout(\storeregister[30][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][4]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[30][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N7
dffeas \storeregister[30][4] (
	.clk(!CLK),
	.d(\storeregister[30][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][4] .is_wysiwyg = "true";
defparam \storeregister[30][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N10
cycloneive_lcell_comb \Mux27~3 (
// Equation(s):
// \Mux27~3_combout  = (temp_imemload_output_23 & ((\Mux27~2_combout  & ((\storeregister[30][4]~q ))) # (!\Mux27~2_combout  & (\storeregister[22][4]~q )))) # (!temp_imemload_output_23 & (\Mux27~2_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux27~2_combout ),
	.datac(\storeregister[22][4]~q ),
	.datad(\storeregister[30][4]~q ),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~3 .lut_mask = 16'hEC64;
defparam \Mux27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N28
cycloneive_lcell_comb \Mux27~6 (
// Equation(s):
// \Mux27~6_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22)))) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & ((\Mux27~3_combout ))) # (!temp_imemload_output_22 & (\Mux27~5_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux27~5_combout ),
	.datac(temp_imemload_output_22),
	.datad(\Mux27~3_combout ),
	.cin(gnd),
	.combout(\Mux27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~6 .lut_mask = 16'hF4A4;
defparam \Mux27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N29
dffeas \storeregister[17][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][4] .is_wysiwyg = "true";
defparam \storeregister[17][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N27
dffeas \storeregister[21][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][4] .is_wysiwyg = "true";
defparam \storeregister[21][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N28
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\storeregister[21][4]~q )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & (\storeregister[17][4]~q )))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[17][4]~q ),
	.datad(\storeregister[21][4]~q ),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hBA98;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N25
dffeas \storeregister[29][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][4] .is_wysiwyg = "true";
defparam \storeregister[29][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N7
dffeas \storeregister[25][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][4] .is_wysiwyg = "true";
defparam \storeregister[25][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N24
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (temp_imemload_output_24 & ((\Mux27~0_combout  & (\storeregister[29][4]~q )) # (!\Mux27~0_combout  & ((\storeregister[25][4]~q ))))) # (!temp_imemload_output_24 & (\Mux27~0_combout ))

	.dataa(temp_imemload_output_24),
	.datab(\Mux27~0_combout ),
	.datac(\storeregister[29][4]~q ),
	.datad(\storeregister[25][4]~q ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hE6C4;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N21
dffeas \storeregister[3][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][4] .is_wysiwyg = "true";
defparam \storeregister[3][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N27
dffeas \storeregister[1][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][4] .is_wysiwyg = "true";
defparam \storeregister[1][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N26
cycloneive_lcell_comb \Mux27~14 (
// Equation(s):
// \Mux27~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[3][4]~q )) # (!temp_imemload_output_22 & ((\storeregister[1][4]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[3][4]~q ),
	.datac(\storeregister[1][4]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux27~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~14 .lut_mask = 16'h88A0;
defparam \Mux27~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N4
cycloneive_lcell_comb \Mux27~15 (
// Equation(s):
// \Mux27~15_combout  = (\Mux27~14_combout ) # ((\storeregister[2][4]~q  & (!temp_imemload_output_21 & temp_imemload_output_22)))

	.dataa(\storeregister[2][4]~q ),
	.datab(temp_imemload_output_21),
	.datac(temp_imemload_output_22),
	.datad(\Mux27~14_combout ),
	.cin(gnd),
	.combout(\Mux27~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~15 .lut_mask = 16'hFF20;
defparam \Mux27~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N2
cycloneive_lcell_comb \storeregister[7][4]~feeder (
// Equation(s):
// \storeregister[7][4]~feeder_combout  = Mux27

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux27),
	.cin(gnd),
	.combout(\storeregister[7][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[7][4]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[7][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N3
dffeas \storeregister[7][4] (
	.clk(!CLK),
	.d(\storeregister[7][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][4] .is_wysiwyg = "true";
defparam \storeregister[7][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y42_N31
dffeas \storeregister[4][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][4] .is_wysiwyg = "true";
defparam \storeregister[4][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y42_N13
dffeas \storeregister[5][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][4] .is_wysiwyg = "true";
defparam \storeregister[5][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N30
cycloneive_lcell_comb \Mux27~12 (
// Equation(s):
// \Mux27~12_combout  = (temp_imemload_output_22 & (temp_imemload_output_21)) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[5][4]~q ))) # (!temp_imemload_output_21 & (\storeregister[4][4]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[4][4]~q ),
	.datad(\storeregister[5][4]~q ),
	.cin(gnd),
	.combout(\Mux27~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~12 .lut_mask = 16'hDC98;
defparam \Mux27~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N24
cycloneive_lcell_comb \Mux27~13 (
// Equation(s):
// \Mux27~13_combout  = (\Mux27~12_combout  & (((\storeregister[7][4]~q ) # (!temp_imemload_output_22)))) # (!\Mux27~12_combout  & (\storeregister[6][4]~q  & ((temp_imemload_output_22))))

	.dataa(\storeregister[6][4]~q ),
	.datab(\storeregister[7][4]~q ),
	.datac(\Mux27~12_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux27~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~13 .lut_mask = 16'hCAF0;
defparam \Mux27~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N18
cycloneive_lcell_comb \Mux27~16 (
// Equation(s):
// \Mux27~16_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\Mux27~13_combout )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & (\Mux27~15_combout )))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\Mux27~15_combout ),
	.datad(\Mux27~13_combout ),
	.cin(gnd),
	.combout(\Mux27~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~16 .lut_mask = 16'hBA98;
defparam \Mux27~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N19
dffeas \storeregister[10][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][4] .is_wysiwyg = "true";
defparam \storeregister[10][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N26
cycloneive_lcell_comb \storeregister[8][4]~feeder (
// Equation(s):
// \storeregister[8][4]~feeder_combout  = Mux27

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux27),
	.cin(gnd),
	.combout(\storeregister[8][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[8][4]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[8][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N27
dffeas \storeregister[8][4] (
	.clk(!CLK),
	.d(\storeregister[8][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][4] .is_wysiwyg = "true";
defparam \storeregister[8][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N18
cycloneive_lcell_comb \Mux27~10 (
// Equation(s):
// \Mux27~10_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[10][4]~q )) # (!temp_imemload_output_22 & ((\storeregister[8][4]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][4]~q ),
	.datad(\storeregister[8][4]~q ),
	.cin(gnd),
	.combout(\Mux27~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~10 .lut_mask = 16'hD9C8;
defparam \Mux27~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N25
dffeas \storeregister[9][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][4] .is_wysiwyg = "true";
defparam \storeregister[9][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N4
cycloneive_lcell_comb \storeregister[11][4]~feeder (
// Equation(s):
// \storeregister[11][4]~feeder_combout  = Mux27

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux27),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[11][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[11][4]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[11][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N5
dffeas \storeregister[11][4] (
	.clk(!CLK),
	.d(\storeregister[11][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][4] .is_wysiwyg = "true";
defparam \storeregister[11][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N24
cycloneive_lcell_comb \Mux27~11 (
// Equation(s):
// \Mux27~11_combout  = (temp_imemload_output_21 & ((\Mux27~10_combout  & ((\storeregister[11][4]~q ))) # (!\Mux27~10_combout  & (\storeregister[9][4]~q )))) # (!temp_imemload_output_21 & (\Mux27~10_combout ))

	.dataa(temp_imemload_output_21),
	.datab(\Mux27~10_combout ),
	.datac(\storeregister[9][4]~q ),
	.datad(\storeregister[11][4]~q ),
	.cin(gnd),
	.combout(\Mux27~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~11 .lut_mask = 16'hEC64;
defparam \Mux27~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N23
dffeas \storeregister[12][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][4] .is_wysiwyg = "true";
defparam \storeregister[12][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N13
dffeas \storeregister[13][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][4] .is_wysiwyg = "true";
defparam \storeregister[13][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N12
cycloneive_lcell_comb \Mux27~17 (
// Equation(s):
// \Mux27~17_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[13][4]~q ))) # (!temp_imemload_output_21 & (\storeregister[12][4]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[12][4]~q ),
	.datac(\storeregister[13][4]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux27~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~17 .lut_mask = 16'hFA44;
defparam \Mux27~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N8
cycloneive_lcell_comb \storeregister[14][4]~feeder (
// Equation(s):
// \storeregister[14][4]~feeder_combout  = Mux27

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux27),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[14][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][4]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[14][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y39_N9
dffeas \storeregister[14][4] (
	.clk(!CLK),
	.d(\storeregister[14][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][4] .is_wysiwyg = "true";
defparam \storeregister[14][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N26
cycloneive_lcell_comb \storeregister[15][4]~feeder (
// Equation(s):
// \storeregister[15][4]~feeder_combout  = Mux27

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux27),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[15][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][4]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[15][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N27
dffeas \storeregister[15][4] (
	.clk(!CLK),
	.d(\storeregister[15][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][4] .is_wysiwyg = "true";
defparam \storeregister[15][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N26
cycloneive_lcell_comb \Mux27~18 (
// Equation(s):
// \Mux27~18_combout  = (\Mux27~17_combout  & (((\storeregister[15][4]~q )) # (!temp_imemload_output_22))) # (!\Mux27~17_combout  & (temp_imemload_output_22 & (\storeregister[14][4]~q )))

	.dataa(\Mux27~17_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[14][4]~q ),
	.datad(\storeregister[15][4]~q ),
	.cin(gnd),
	.combout(\Mux27~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~18 .lut_mask = 16'hEA62;
defparam \Mux27~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N25
dffeas \storeregister[20][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][3] .is_wysiwyg = "true";
defparam \storeregister[20][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N19
dffeas \storeregister[16][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][3] .is_wysiwyg = "true";
defparam \storeregister[16][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N24
cycloneive_lcell_comb \Mux28~4 (
// Equation(s):
// \Mux28~4_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\storeregister[20][3]~q )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & ((\storeregister[16][3]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[20][3]~q ),
	.datad(\storeregister[16][3]~q ),
	.cin(gnd),
	.combout(\Mux28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~4 .lut_mask = 16'hB9A8;
defparam \Mux28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N30
cycloneive_lcell_comb \storeregister[28][3]~feeder (
// Equation(s):
// \storeregister[28][3]~feeder_combout  = Mux28

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux28),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[28][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][3]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[28][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N31
dffeas \storeregister[28][3] (
	.clk(!CLK),
	.d(\storeregister[28][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][3] .is_wysiwyg = "true";
defparam \storeregister[28][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N8
cycloneive_lcell_comb \Mux28~5 (
// Equation(s):
// \Mux28~5_combout  = (\Mux28~4_combout  & (((\storeregister[28][3]~q ) # (!temp_imemload_output_24)))) # (!\Mux28~4_combout  & (\storeregister[24][3]~q  & ((temp_imemload_output_24))))

	.dataa(\storeregister[24][3]~q ),
	.datab(\Mux28~4_combout ),
	.datac(\storeregister[28][3]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~5 .lut_mask = 16'hE2CC;
defparam \Mux28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N16
cycloneive_lcell_comb \storeregister[22][3]~feeder (
// Equation(s):
// \storeregister[22][3]~feeder_combout  = Mux28

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux28),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[22][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[22][3]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[22][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N17
dffeas \storeregister[22][3] (
	.clk(!CLK),
	.d(\storeregister[22][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][3] .is_wysiwyg = "true";
defparam \storeregister[22][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N19
dffeas \storeregister[18][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][3] .is_wysiwyg = "true";
defparam \storeregister[18][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N18
cycloneive_lcell_comb \Mux28~2 (
// Equation(s):
// \Mux28~2_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[22][3]~q )) # (!temp_imemload_output_23 & ((\storeregister[18][3]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[22][3]~q ),
	.datac(\storeregister[18][3]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~2 .lut_mask = 16'hEE50;
defparam \Mux28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N17
dffeas \storeregister[26][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][3] .is_wysiwyg = "true";
defparam \storeregister[26][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N10
cycloneive_lcell_comb \Mux28~3 (
// Equation(s):
// \Mux28~3_combout  = (temp_imemload_output_24 & ((\Mux28~2_combout  & (\storeregister[30][3]~q )) # (!\Mux28~2_combout  & ((\storeregister[26][3]~q ))))) # (!temp_imemload_output_24 & (((\Mux28~2_combout ))))

	.dataa(\storeregister[30][3]~q ),
	.datab(temp_imemload_output_24),
	.datac(\Mux28~2_combout ),
	.datad(\storeregister[26][3]~q ),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~3 .lut_mask = 16'hBCB0;
defparam \Mux28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N14
cycloneive_lcell_comb \Mux28~6 (
// Equation(s):
// \Mux28~6_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21) # (\Mux28~3_combout )))) # (!temp_imemload_output_22 & (\Mux28~5_combout  & (!temp_imemload_output_21)))

	.dataa(\Mux28~5_combout ),
	.datab(temp_imemload_output_22),
	.datac(temp_imemload_output_21),
	.datad(\Mux28~3_combout ),
	.cin(gnd),
	.combout(\Mux28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~6 .lut_mask = 16'hCEC2;
defparam \Mux28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N0
cycloneive_lcell_comb \storeregister[25][3]~feeder (
// Equation(s):
// \storeregister[25][3]~feeder_combout  = Mux28

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux28),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[25][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[25][3]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[25][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N1
dffeas \storeregister[25][3] (
	.clk(!CLK),
	.d(\storeregister[25][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][3] .is_wysiwyg = "true";
defparam \storeregister[25][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N7
dffeas \storeregister[17][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][3] .is_wysiwyg = "true";
defparam \storeregister[17][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N6
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (temp_imemload_output_24 & ((\storeregister[25][3]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[17][3]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[25][3]~q ),
	.datac(\storeregister[17][3]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hAAD8;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N29
dffeas \storeregister[29][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][3] .is_wysiwyg = "true";
defparam \storeregister[29][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N29
dffeas \storeregister[21][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][3] .is_wysiwyg = "true";
defparam \storeregister[21][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N28
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (\Mux28~0_combout  & (((\storeregister[29][3]~q )) # (!temp_imemload_output_23))) # (!\Mux28~0_combout  & (temp_imemload_output_23 & ((\storeregister[21][3]~q ))))

	.dataa(\Mux28~0_combout ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[29][3]~q ),
	.datad(\storeregister[21][3]~q ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hE6A2;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N26
cycloneive_lcell_comb \storeregister[27][3]~feeder (
// Equation(s):
// \storeregister[27][3]~feeder_combout  = Mux28

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux28),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][3]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N27
dffeas \storeregister[27][3] (
	.clk(!CLK),
	.d(\storeregister[27][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][3] .is_wysiwyg = "true";
defparam \storeregister[27][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N20
cycloneive_lcell_comb \Mux28~7 (
// Equation(s):
// \Mux28~7_combout  = (temp_imemload_output_24 & (((\storeregister[27][3]~q ) # (temp_imemload_output_23)))) # (!temp_imemload_output_24 & (\storeregister[19][3]~q  & ((!temp_imemload_output_23))))

	.dataa(\storeregister[19][3]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[27][3]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~7 .lut_mask = 16'hCCE2;
defparam \Mux28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N19
dffeas \storeregister[23][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][3] .is_wysiwyg = "true";
defparam \storeregister[23][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N2
cycloneive_lcell_comb \storeregister[31][3]~feeder (
// Equation(s):
// \storeregister[31][3]~feeder_combout  = Mux28

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux28),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[31][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][3]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[31][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N3
dffeas \storeregister[31][3] (
	.clk(!CLK),
	.d(\storeregister[31][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][3] .is_wysiwyg = "true";
defparam \storeregister[31][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N18
cycloneive_lcell_comb \Mux28~8 (
// Equation(s):
// \Mux28~8_combout  = (\Mux28~7_combout  & (((\storeregister[31][3]~q )) # (!temp_imemload_output_23))) # (!\Mux28~7_combout  & (temp_imemload_output_23 & (\storeregister[23][3]~q )))

	.dataa(\Mux28~7_combout ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[23][3]~q ),
	.datad(\storeregister[31][3]~q ),
	.cin(gnd),
	.combout(\Mux28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~8 .lut_mask = 16'hEA62;
defparam \Mux28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N6
cycloneive_lcell_comb \storeregister[6][3]~feeder (
// Equation(s):
// \storeregister[6][3]~feeder_combout  = Mux28

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux28),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[6][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[6][3]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[6][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N7
dffeas \storeregister[6][3] (
	.clk(!CLK),
	.d(\storeregister[6][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][3] .is_wysiwyg = "true";
defparam \storeregister[6][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y42_N1
dffeas \storeregister[5][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][3] .is_wysiwyg = "true";
defparam \storeregister[5][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y42_N11
dffeas \storeregister[4][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][3] .is_wysiwyg = "true";
defparam \storeregister[4][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N0
cycloneive_lcell_comb \Mux28~10 (
// Equation(s):
// \Mux28~10_combout  = (temp_imemload_output_22 & (temp_imemload_output_21)) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & (\storeregister[5][3]~q )) # (!temp_imemload_output_21 & ((\storeregister[4][3]~q )))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[5][3]~q ),
	.datad(\storeregister[4][3]~q ),
	.cin(gnd),
	.combout(\Mux28~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~10 .lut_mask = 16'hD9C8;
defparam \Mux28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N10
cycloneive_lcell_comb \storeregister[7][3]~feeder (
// Equation(s):
// \storeregister[7][3]~feeder_combout  = Mux28

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux28),
	.cin(gnd),
	.combout(\storeregister[7][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[7][3]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[7][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N11
dffeas \storeregister[7][3] (
	.clk(!CLK),
	.d(\storeregister[7][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][3] .is_wysiwyg = "true";
defparam \storeregister[7][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N12
cycloneive_lcell_comb \Mux28~11 (
// Equation(s):
// \Mux28~11_combout  = (temp_imemload_output_22 & ((\Mux28~10_combout  & ((\storeregister[7][3]~q ))) # (!\Mux28~10_combout  & (\storeregister[6][3]~q )))) # (!temp_imemload_output_22 & (((\Mux28~10_combout ))))

	.dataa(\storeregister[6][3]~q ),
	.datab(temp_imemload_output_22),
	.datac(\Mux28~10_combout ),
	.datad(\storeregister[7][3]~q ),
	.cin(gnd),
	.combout(\Mux28~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~11 .lut_mask = 16'hF838;
defparam \Mux28~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N24
cycloneive_lcell_comb \storeregister[9][3]~feeder (
// Equation(s):
// \storeregister[9][3]~feeder_combout  = Mux28

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux28),
	.cin(gnd),
	.combout(\storeregister[9][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[9][3]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[9][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N25
dffeas \storeregister[9][3] (
	.clk(!CLK),
	.d(\storeregister[9][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][3] .is_wysiwyg = "true";
defparam \storeregister[9][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N1
dffeas \storeregister[11][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][3] .is_wysiwyg = "true";
defparam \storeregister[11][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N5
dffeas \storeregister[10][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][3] .is_wysiwyg = "true";
defparam \storeregister[10][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N7
dffeas \storeregister[8][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][3] .is_wysiwyg = "true";
defparam \storeregister[8][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N6
cycloneive_lcell_comb \Mux28~12 (
// Equation(s):
// \Mux28~12_combout  = (temp_imemload_output_22 & ((\storeregister[10][3]~q ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((\storeregister[8][3]~q  & !temp_imemload_output_21))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[10][3]~q ),
	.datac(\storeregister[8][3]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux28~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~12 .lut_mask = 16'hAAD8;
defparam \Mux28~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N0
cycloneive_lcell_comb \Mux28~13 (
// Equation(s):
// \Mux28~13_combout  = (temp_imemload_output_21 & ((\Mux28~12_combout  & ((\storeregister[11][3]~q ))) # (!\Mux28~12_combout  & (\storeregister[9][3]~q )))) # (!temp_imemload_output_21 & (((\Mux28~12_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[9][3]~q ),
	.datac(\storeregister[11][3]~q ),
	.datad(\Mux28~12_combout ),
	.cin(gnd),
	.combout(\Mux28~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~13 .lut_mask = 16'hF588;
defparam \Mux28~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N31
dffeas \storeregister[2][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][3] .is_wysiwyg = "true";
defparam \storeregister[2][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N24
cycloneive_lcell_comb \Mux28~15 (
// Equation(s):
// \Mux28~15_combout  = (\Mux28~14_combout ) # ((temp_imemload_output_22 & (\storeregister[2][3]~q  & !temp_imemload_output_21)))

	.dataa(\Mux28~14_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][3]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux28~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~15 .lut_mask = 16'hAAEA;
defparam \Mux28~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N26
cycloneive_lcell_comb \Mux28~16 (
// Equation(s):
// \Mux28~16_combout  = (temp_imemload_output_24 & ((temp_imemload_output_23) # ((\Mux28~13_combout )))) # (!temp_imemload_output_24 & (!temp_imemload_output_23 & ((\Mux28~15_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\Mux28~13_combout ),
	.datad(\Mux28~15_combout ),
	.cin(gnd),
	.combout(\Mux28~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~16 .lut_mask = 16'hB9A8;
defparam \Mux28~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N17
dffeas \storeregister[15][3] (
	.clk(!CLK),
	.d(Mux28),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][3] .is_wysiwyg = "true";
defparam \storeregister[15][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y42_N13
dffeas \storeregister[14][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][3] .is_wysiwyg = "true";
defparam \storeregister[14][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N15
dffeas \storeregister[12][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][3] .is_wysiwyg = "true";
defparam \storeregister[12][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N21
dffeas \storeregister[13][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][3] .is_wysiwyg = "true";
defparam \storeregister[13][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N20
cycloneive_lcell_comb \Mux28~17 (
// Equation(s):
// \Mux28~17_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[13][3]~q ))) # (!temp_imemload_output_21 & (\storeregister[12][3]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[12][3]~q ),
	.datac(\storeregister[13][3]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux28~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~17 .lut_mask = 16'hFA44;
defparam \Mux28~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N12
cycloneive_lcell_comb \Mux28~18 (
// Equation(s):
// \Mux28~18_combout  = (temp_imemload_output_22 & ((\Mux28~17_combout  & (\storeregister[15][3]~q )) # (!\Mux28~17_combout  & ((\storeregister[14][3]~q ))))) # (!temp_imemload_output_22 & (((\Mux28~17_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[15][3]~q ),
	.datac(\storeregister[14][3]~q ),
	.datad(\Mux28~17_combout ),
	.cin(gnd),
	.combout(\Mux28~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~18 .lut_mask = 16'hDDA0;
defparam \Mux28~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N0
cycloneive_lcell_comb \Mux61~4 (
// Equation(s):
// \Mux61~4_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\storeregister[20][2]~q )) # (!temp_imemload_output_18 & ((\storeregister[16][2]~q )))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[20][2]~q ),
	.datad(\storeregister[16][2]~q ),
	.cin(gnd),
	.combout(\Mux61~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~4 .lut_mask = 16'hD9C8;
defparam \Mux61~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N0
cycloneive_lcell_comb \Mux61~5 (
// Equation(s):
// \Mux61~5_combout  = (\Mux61~4_combout  & ((\storeregister[28][2]~q ) # ((!temp_imemload_output_19)))) # (!\Mux61~4_combout  & (((temp_imemload_output_19 & \storeregister[24][2]~q ))))

	.dataa(\storeregister[28][2]~q ),
	.datab(\Mux61~4_combout ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[24][2]~q ),
	.cin(gnd),
	.combout(\Mux61~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~5 .lut_mask = 16'hBC8C;
defparam \Mux61~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N7
dffeas \storeregister[22][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][2] .is_wysiwyg = "true";
defparam \storeregister[22][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N6
cycloneive_lcell_comb \Mux61~2 (
// Equation(s):
// \Mux61~2_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[22][2]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[18][2]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[22][2]~q ),
	.datad(\storeregister[18][2]~q ),
	.cin(gnd),
	.combout(\Mux61~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~2 .lut_mask = 16'hB9A8;
defparam \Mux61~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N30
cycloneive_lcell_comb \Mux61~3 (
// Equation(s):
// \Mux61~3_combout  = (temp_imemload_output_19 & ((\Mux61~2_combout  & (\storeregister[30][2]~q )) # (!\Mux61~2_combout  & ((\storeregister[26][2]~q ))))) # (!temp_imemload_output_19 & (((\Mux61~2_combout ))))

	.dataa(\storeregister[30][2]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[26][2]~q ),
	.datad(\Mux61~2_combout ),
	.cin(gnd),
	.combout(\Mux61~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~3 .lut_mask = 16'hBBC0;
defparam \Mux61~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N12
cycloneive_lcell_comb \Mux61~6 (
// Equation(s):
// \Mux61~6_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16) # (\Mux61~3_combout )))) # (!temp_imemload_output_17 & (\Mux61~5_combout  & (!temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux61~5_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux61~3_combout ),
	.cin(gnd),
	.combout(\Mux61~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~6 .lut_mask = 16'hAEA4;
defparam \Mux61~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N21
dffeas \storeregister[21][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][2] .is_wysiwyg = "true";
defparam \storeregister[21][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N2
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (temp_imemload_output_19 & (((\storeregister[25][2]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[17][2]~q  & ((!temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[17][2]~q ),
	.datac(\storeregister[25][2]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'hAAE4;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N20
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (temp_imemload_output_18 & ((\Mux61~0_combout  & (\storeregister[29][2]~q )) # (!\Mux61~0_combout  & ((\storeregister[21][2]~q ))))) # (!temp_imemload_output_18 & (((\Mux61~0_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[29][2]~q ),
	.datac(\storeregister[21][2]~q ),
	.datad(\Mux61~0_combout ),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hDDA0;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N4
cycloneive_lcell_comb \Mux61~7 (
// Equation(s):
// \Mux61~7_combout  = (temp_imemload_output_19 & ((\storeregister[27][2]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\storeregister[19][2]~q  & !temp_imemload_output_18))))

	.dataa(\storeregister[27][2]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[19][2]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux61~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~7 .lut_mask = 16'hCCB8;
defparam \Mux61~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N28
cycloneive_lcell_comb \Mux61~8 (
// Equation(s):
// \Mux61~8_combout  = (temp_imemload_output_18 & ((\Mux61~7_combout  & (\storeregister[31][2]~q )) # (!\Mux61~7_combout  & ((\storeregister[23][2]~q ))))) # (!temp_imemload_output_18 & (\Mux61~7_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux61~7_combout ),
	.datac(\storeregister[31][2]~q ),
	.datad(\storeregister[23][2]~q ),
	.cin(gnd),
	.combout(\Mux61~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~8 .lut_mask = 16'hE6C4;
defparam \Mux61~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N4
cycloneive_lcell_comb \Mux61~14 (
// Equation(s):
// \Mux61~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][2]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][2]~q )))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[3][2]~q ),
	.datad(\storeregister[1][2]~q ),
	.cin(gnd),
	.combout(\Mux61~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~14 .lut_mask = 16'hA280;
defparam \Mux61~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N10
cycloneive_lcell_comb \storeregister[2][2]~feeder (
// Equation(s):
// \storeregister[2][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux29),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[2][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[2][2]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[2][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N11
dffeas \storeregister[2][2] (
	.clk(!CLK),
	.d(\storeregister[2][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][2] .is_wysiwyg = "true";
defparam \storeregister[2][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N6
cycloneive_lcell_comb \Mux61~15 (
// Equation(s):
// \Mux61~15_combout  = (\Mux61~14_combout ) # ((!temp_imemload_output_16 & (temp_imemload_output_17 & \storeregister[2][2]~q )))

	.dataa(temp_imemload_output_16),
	.datab(\Mux61~14_combout ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[2][2]~q ),
	.cin(gnd),
	.combout(\Mux61~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~15 .lut_mask = 16'hDCCC;
defparam \Mux61~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N20
cycloneive_lcell_comb \Mux61~12 (
// Equation(s):
// \Mux61~12_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[10][2]~q ))) # (!temp_imemload_output_17 & (\storeregister[8][2]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[8][2]~q ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[10][2]~q ),
	.cin(gnd),
	.combout(\Mux61~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~12 .lut_mask = 16'hF4A4;
defparam \Mux61~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N8
cycloneive_lcell_comb \Mux61~13 (
// Equation(s):
// \Mux61~13_combout  = (temp_imemload_output_16 & ((\Mux61~12_combout  & ((\storeregister[11][2]~q ))) # (!\Mux61~12_combout  & (\storeregister[9][2]~q )))) # (!temp_imemload_output_16 & (\Mux61~12_combout ))

	.dataa(temp_imemload_output_16),
	.datab(\Mux61~12_combout ),
	.datac(\storeregister[9][2]~q ),
	.datad(\storeregister[11][2]~q ),
	.cin(gnd),
	.combout(\Mux61~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~13 .lut_mask = 16'hEC64;
defparam \Mux61~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N20
cycloneive_lcell_comb \Mux61~16 (
// Equation(s):
// \Mux61~16_combout  = (temp_imemload_output_19 & (((\Mux61~13_combout ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\Mux61~15_combout  & ((!temp_imemload_output_18))))

	.dataa(\Mux61~15_combout ),
	.datab(\Mux61~13_combout ),
	.datac(temp_imemload_output_19),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux61~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~16 .lut_mask = 16'hF0CA;
defparam \Mux61~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N30
cycloneive_lcell_comb \storeregister[7][2]~feeder (
// Equation(s):
// \storeregister[7][2]~feeder_combout  = Mux29

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux29),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[7][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[7][2]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[7][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N31
dffeas \storeregister[7][2] (
	.clk(!CLK),
	.d(\storeregister[7][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][2] .is_wysiwyg = "true";
defparam \storeregister[7][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N28
cycloneive_lcell_comb \Mux61~10 (
// Equation(s):
// \Mux61~10_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[5][2]~q ))) # (!temp_imemload_output_16 & (\storeregister[4][2]~q ))))

	.dataa(\storeregister[4][2]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][2]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux61~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~10 .lut_mask = 16'hFC22;
defparam \Mux61~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N14
cycloneive_lcell_comb \Mux61~11 (
// Equation(s):
// \Mux61~11_combout  = (temp_imemload_output_17 & ((\Mux61~10_combout  & ((\storeregister[7][2]~q ))) # (!\Mux61~10_combout  & (\storeregister[6][2]~q )))) # (!temp_imemload_output_17 & (((\Mux61~10_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[6][2]~q ),
	.datac(\storeregister[7][2]~q ),
	.datad(\Mux61~10_combout ),
	.cin(gnd),
	.combout(\Mux61~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~11 .lut_mask = 16'hF588;
defparam \Mux61~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N2
cycloneive_lcell_comb \Mux61~17 (
// Equation(s):
// \Mux61~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][2]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][2]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[12][2]~q ),
	.datad(\storeregister[13][2]~q ),
	.cin(gnd),
	.combout(\Mux61~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~17 .lut_mask = 16'hDC98;
defparam \Mux61~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N6
cycloneive_lcell_comb \Mux61~18 (
// Equation(s):
// \Mux61~18_combout  = (temp_imemload_output_17 & ((\Mux61~17_combout  & (\storeregister[15][2]~q )) # (!\Mux61~17_combout  & ((\storeregister[14][2]~q ))))) # (!temp_imemload_output_17 & (((\Mux61~17_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[15][2]~q ),
	.datac(\Mux61~17_combout ),
	.datad(\storeregister[14][2]~q ),
	.cin(gnd),
	.combout(\Mux61~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~18 .lut_mask = 16'hDAD0;
defparam \Mux61~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N3
dffeas \storeregister[23][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][8] .is_wysiwyg = "true";
defparam \storeregister[23][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N9
dffeas \storeregister[19][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][8] .is_wysiwyg = "true";
defparam \storeregister[19][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N2
cycloneive_lcell_comb \Mux23~7 (
// Equation(s):
// \Mux23~7_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[23][8]~q )) # (!temp_imemload_output_23 & ((\storeregister[19][8]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[23][8]~q ),
	.datad(\storeregister[19][8]~q ),
	.cin(gnd),
	.combout(\Mux23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~7 .lut_mask = 16'hD9C8;
defparam \Mux23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N8
cycloneive_lcell_comb \storeregister[27][8]~feeder (
// Equation(s):
// \storeregister[27][8]~feeder_combout  = Mux23

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux23),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][8]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N9
dffeas \storeregister[27][8] (
	.clk(!CLK),
	.d(\storeregister[27][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][8] .is_wysiwyg = "true";
defparam \storeregister[27][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N18
cycloneive_lcell_comb \storeregister[31][8]~feeder (
// Equation(s):
// \storeregister[31][8]~feeder_combout  = Mux23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux23),
	.cin(gnd),
	.combout(\storeregister[31][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][8]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[31][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N19
dffeas \storeregister[31][8] (
	.clk(!CLK),
	.d(\storeregister[31][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][8] .is_wysiwyg = "true";
defparam \storeregister[31][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N20
cycloneive_lcell_comb \Mux23~8 (
// Equation(s):
// \Mux23~8_combout  = (\Mux23~7_combout  & (((\storeregister[31][8]~q )) # (!temp_imemload_output_24))) # (!\Mux23~7_combout  & (temp_imemload_output_24 & (\storeregister[27][8]~q )))

	.dataa(\Mux23~7_combout ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[27][8]~q ),
	.datad(\storeregister[31][8]~q ),
	.cin(gnd),
	.combout(\Mux23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~8 .lut_mask = 16'hEA62;
defparam \Mux23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N17
dffeas \storeregister[26][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][8] .is_wysiwyg = "true";
defparam \storeregister[26][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N0
cycloneive_lcell_comb \storeregister[18][8]~feeder (
// Equation(s):
// \storeregister[18][8]~feeder_combout  = Mux23

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux23),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[18][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[18][8]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[18][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N1
dffeas \storeregister[18][8] (
	.clk(!CLK),
	.d(\storeregister[18][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][8] .is_wysiwyg = "true";
defparam \storeregister[18][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N6
cycloneive_lcell_comb \Mux23~2 (
// Equation(s):
// \Mux23~2_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[26][8]~q )) # (!temp_imemload_output_24 & ((\storeregister[18][8]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[26][8]~q ),
	.datad(\storeregister[18][8]~q ),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~2 .lut_mask = 16'hD9C8;
defparam \Mux23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N16
cycloneive_lcell_comb \storeregister[30][8]~feeder (
// Equation(s):
// \storeregister[30][8]~feeder_combout  = Mux23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux23),
	.cin(gnd),
	.combout(\storeregister[30][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][8]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[30][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N17
dffeas \storeregister[30][8] (
	.clk(!CLK),
	.d(\storeregister[30][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][8] .is_wysiwyg = "true";
defparam \storeregister[30][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N26
cycloneive_lcell_comb \Mux23~3 (
// Equation(s):
// \Mux23~3_combout  = (temp_imemload_output_23 & ((\Mux23~2_combout  & ((\storeregister[30][8]~q ))) # (!\Mux23~2_combout  & (\storeregister[22][8]~q )))) # (!temp_imemload_output_23 & (((\Mux23~2_combout ))))

	.dataa(\storeregister[22][8]~q ),
	.datab(temp_imemload_output_23),
	.datac(\Mux23~2_combout ),
	.datad(\storeregister[30][8]~q ),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~3 .lut_mask = 16'hF838;
defparam \Mux23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N14
cycloneive_lcell_comb \storeregister[28][8]~feeder (
// Equation(s):
// \storeregister[28][8]~feeder_combout  = Mux23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux23),
	.cin(gnd),
	.combout(\storeregister[28][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][8]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[28][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N15
dffeas \storeregister[28][8] (
	.clk(!CLK),
	.d(\storeregister[28][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][8] .is_wysiwyg = "true";
defparam \storeregister[28][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N28
cycloneive_lcell_comb \storeregister[20][8]~feeder (
// Equation(s):
// \storeregister[20][8]~feeder_combout  = Mux23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux23),
	.cin(gnd),
	.combout(\storeregister[20][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][8]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[20][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N29
dffeas \storeregister[20][8] (
	.clk(!CLK),
	.d(\storeregister[20][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][8] .is_wysiwyg = "true";
defparam \storeregister[20][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N12
cycloneive_lcell_comb \Mux23~5 (
// Equation(s):
// \Mux23~5_combout  = (\Mux23~4_combout  & (((\storeregister[28][8]~q )) # (!temp_imemload_output_23))) # (!\Mux23~4_combout  & (temp_imemload_output_23 & ((\storeregister[20][8]~q ))))

	.dataa(\Mux23~4_combout ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[28][8]~q ),
	.datad(\storeregister[20][8]~q ),
	.cin(gnd),
	.combout(\Mux23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~5 .lut_mask = 16'hE6A2;
defparam \Mux23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N22
cycloneive_lcell_comb \Mux23~6 (
// Equation(s):
// \Mux23~6_combout  = (temp_imemload_output_22 & ((\Mux23~3_combout ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((!temp_imemload_output_21 & \Mux23~5_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(\Mux23~3_combout ),
	.datac(temp_imemload_output_21),
	.datad(\Mux23~5_combout ),
	.cin(gnd),
	.combout(\Mux23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~6 .lut_mask = 16'hADA8;
defparam \Mux23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N4
cycloneive_lcell_comb \storeregister[21][8]~feeder (
// Equation(s):
// \storeregister[21][8]~feeder_combout  = Mux23

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux23),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[21][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][8]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[21][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N5
dffeas \storeregister[21][8] (
	.clk(!CLK),
	.d(\storeregister[21][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][8] .is_wysiwyg = "true";
defparam \storeregister[21][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N0
cycloneive_lcell_comb \storeregister[17][8]~feeder (
// Equation(s):
// \storeregister[17][8]~feeder_combout  = Mux23

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux23),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[17][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[17][8]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[17][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N1
dffeas \storeregister[17][8] (
	.clk(!CLK),
	.d(\storeregister[17][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][8] .is_wysiwyg = "true";
defparam \storeregister[17][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N6
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[21][8]~q )) # (!temp_imemload_output_23 & ((\storeregister[17][8]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[21][8]~q ),
	.datac(temp_imemload_output_23),
	.datad(\storeregister[17][8]~q ),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hE5E0;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N7
dffeas \storeregister[25][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][8] .is_wysiwyg = "true";
defparam \storeregister[25][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N30
cycloneive_lcell_comb \storeregister[29][8]~feeder (
// Equation(s):
// \storeregister[29][8]~feeder_combout  = Mux23

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux23),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[29][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][8]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[29][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y37_N31
dffeas \storeregister[29][8] (
	.clk(!CLK),
	.d(\storeregister[29][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][8] .is_wysiwyg = "true";
defparam \storeregister[29][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N6
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (\Mux23~0_combout  & (((\storeregister[29][8]~q )) # (!temp_imemload_output_24))) # (!\Mux23~0_combout  & (temp_imemload_output_24 & (\storeregister[25][8]~q )))

	.dataa(\Mux23~0_combout ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[25][8]~q ),
	.datad(\storeregister[29][8]~q ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hEA62;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N7
dffeas \storeregister[11][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][8] .is_wysiwyg = "true";
defparam \storeregister[11][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N27
dffeas \storeregister[9][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][8] .is_wysiwyg = "true";
defparam \storeregister[9][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N5
dffeas \storeregister[8][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][8] .is_wysiwyg = "true";
defparam \storeregister[8][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N5
dffeas \storeregister[10][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][8] .is_wysiwyg = "true";
defparam \storeregister[10][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N4
cycloneive_lcell_comb \Mux23~10 (
// Equation(s):
// \Mux23~10_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22)))) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[10][8]~q ))) # (!temp_imemload_output_22 & (\storeregister[8][8]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[8][8]~q ),
	.datac(\storeregister[10][8]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux23~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~10 .lut_mask = 16'hFA44;
defparam \Mux23~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N26
cycloneive_lcell_comb \Mux23~11 (
// Equation(s):
// \Mux23~11_combout  = (temp_imemload_output_21 & ((\Mux23~10_combout  & (\storeregister[11][8]~q )) # (!\Mux23~10_combout  & ((\storeregister[9][8]~q ))))) # (!temp_imemload_output_21 & (((\Mux23~10_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[11][8]~q ),
	.datac(\storeregister[9][8]~q ),
	.datad(\Mux23~10_combout ),
	.cin(gnd),
	.combout(\Mux23~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~11 .lut_mask = 16'hDDA0;
defparam \Mux23~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N17
dffeas \storeregister[7][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][8] .is_wysiwyg = "true";
defparam \storeregister[7][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y42_N29
dffeas \storeregister[6][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][8] .is_wysiwyg = "true";
defparam \storeregister[6][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N16
cycloneive_lcell_comb \Mux23~13 (
// Equation(s):
// \Mux23~13_combout  = (\Mux23~12_combout  & (((\storeregister[7][8]~q )) # (!temp_imemload_output_22))) # (!\Mux23~12_combout  & (temp_imemload_output_22 & ((\storeregister[6][8]~q ))))

	.dataa(\Mux23~12_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[7][8]~q ),
	.datad(\storeregister[6][8]~q ),
	.cin(gnd),
	.combout(\Mux23~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~13 .lut_mask = 16'hE6A2;
defparam \Mux23~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N11
dffeas \storeregister[2][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][8] .is_wysiwyg = "true";
defparam \storeregister[2][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N24
cycloneive_lcell_comb \Mux23~15 (
// Equation(s):
// \Mux23~15_combout  = (\Mux23~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][8]~q )))

	.dataa(\Mux23~14_combout ),
	.datab(temp_imemload_output_21),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[2][8]~q ),
	.cin(gnd),
	.combout(\Mux23~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~15 .lut_mask = 16'hBAAA;
defparam \Mux23~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N14
cycloneive_lcell_comb \Mux23~16 (
// Equation(s):
// \Mux23~16_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\Mux23~13_combout )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & ((\Mux23~15_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\Mux23~13_combout ),
	.datad(\Mux23~15_combout ),
	.cin(gnd),
	.combout(\Mux23~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~16 .lut_mask = 16'hB9A8;
defparam \Mux23~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N10
cycloneive_lcell_comb \storeregister[14][8]~feeder (
// Equation(s):
// \storeregister[14][8]~feeder_combout  = Mux23

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux23),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[14][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][8]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[14][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y40_N11
dffeas \storeregister[14][8] (
	.clk(!CLK),
	.d(\storeregister[14][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][8] .is_wysiwyg = "true";
defparam \storeregister[14][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N5
dffeas \storeregister[12][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][8] .is_wysiwyg = "true";
defparam \storeregister[12][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N23
dffeas \storeregister[13][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][8] .is_wysiwyg = "true";
defparam \storeregister[13][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N22
cycloneive_lcell_comb \Mux23~17 (
// Equation(s):
// \Mux23~17_combout  = (temp_imemload_output_21 & (((\storeregister[13][8]~q ) # (temp_imemload_output_22)))) # (!temp_imemload_output_21 & (\storeregister[12][8]~q  & ((!temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[12][8]~q ),
	.datac(\storeregister[13][8]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux23~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~17 .lut_mask = 16'hAAE4;
defparam \Mux23~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y40_N21
dffeas \storeregister[15][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][8] .is_wysiwyg = "true";
defparam \storeregister[15][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N6
cycloneive_lcell_comb \Mux23~18 (
// Equation(s):
// \Mux23~18_combout  = (\Mux23~17_combout  & (((\storeregister[15][8]~q ) # (!temp_imemload_output_22)))) # (!\Mux23~17_combout  & (\storeregister[14][8]~q  & (temp_imemload_output_22)))

	.dataa(\storeregister[14][8]~q ),
	.datab(\Mux23~17_combout ),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[15][8]~q ),
	.cin(gnd),
	.combout(\Mux23~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~18 .lut_mask = 16'hEC2C;
defparam \Mux23~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N31
dffeas \storeregister[25][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][7] .is_wysiwyg = "true";
defparam \storeregister[25][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N18
cycloneive_lcell_comb \storeregister[17][7]~feeder (
// Equation(s):
// \storeregister[17][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux24),
	.cin(gnd),
	.combout(\storeregister[17][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[17][7]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[17][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N19
dffeas \storeregister[17][7] (
	.clk(!CLK),
	.d(\storeregister[17][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][7] .is_wysiwyg = "true";
defparam \storeregister[17][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N30
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[25][7]~q )) # (!temp_imemload_output_24 & ((\storeregister[17][7]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[25][7]~q ),
	.datad(\storeregister[17][7]~q ),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hD9C8;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N16
cycloneive_lcell_comb \storeregister[29][7]~feeder (
// Equation(s):
// \storeregister[29][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux24),
	.cin(gnd),
	.combout(\storeregister[29][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][7]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[29][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N17
dffeas \storeregister[29][7] (
	.clk(!CLK),
	.d(\storeregister[29][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][7] .is_wysiwyg = "true";
defparam \storeregister[29][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N12
cycloneive_lcell_comb \storeregister[21][7]~feeder (
// Equation(s):
// \storeregister[21][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux24),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[21][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][7]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[21][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N13
dffeas \storeregister[21][7] (
	.clk(!CLK),
	.d(\storeregister[21][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][7] .is_wysiwyg = "true";
defparam \storeregister[21][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N6
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (temp_imemload_output_23 & ((\Mux24~0_combout  & (\storeregister[29][7]~q )) # (!\Mux24~0_combout  & ((\storeregister[21][7]~q ))))) # (!temp_imemload_output_23 & (\Mux24~0_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux24~0_combout ),
	.datac(\storeregister[29][7]~q ),
	.datad(\storeregister[21][7]~q ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hE6C4;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N20
cycloneive_lcell_comb \storeregister[23][7]~feeder (
// Equation(s):
// \storeregister[23][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux24),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[23][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][7]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[23][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N21
dffeas \storeregister[23][7] (
	.clk(!CLK),
	.d(\storeregister[23][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][7] .is_wysiwyg = "true";
defparam \storeregister[23][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N0
cycloneive_lcell_comb \storeregister[27][7]~feeder (
// Equation(s):
// \storeregister[27][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux24),
	.cin(gnd),
	.combout(\storeregister[27][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][7]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[27][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N1
dffeas \storeregister[27][7] (
	.clk(!CLK),
	.d(\storeregister[27][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][7] .is_wysiwyg = "true";
defparam \storeregister[27][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N3
dffeas \storeregister[19][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][7] .is_wysiwyg = "true";
defparam \storeregister[19][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N2
cycloneive_lcell_comb \Mux24~7 (
// Equation(s):
// \Mux24~7_combout  = (temp_imemload_output_24 & ((\storeregister[27][7]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((!temp_imemload_output_23 & \storeregister[19][7]~q ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[27][7]~q ),
	.datac(temp_imemload_output_23),
	.datad(\storeregister[19][7]~q ),
	.cin(gnd),
	.combout(\Mux24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~7 .lut_mask = 16'hADA8;
defparam \Mux24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N4
cycloneive_lcell_comb \storeregister[31][7]~feeder (
// Equation(s):
// \storeregister[31][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux24),
	.cin(gnd),
	.combout(\storeregister[31][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][7]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[31][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N5
dffeas \storeregister[31][7] (
	.clk(!CLK),
	.d(\storeregister[31][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][7] .is_wysiwyg = "true";
defparam \storeregister[31][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N26
cycloneive_lcell_comb \Mux24~8 (
// Equation(s):
// \Mux24~8_combout  = (\Mux24~7_combout  & (((\storeregister[31][7]~q ) # (!temp_imemload_output_23)))) # (!\Mux24~7_combout  & (\storeregister[23][7]~q  & ((temp_imemload_output_23))))

	.dataa(\storeregister[23][7]~q ),
	.datab(\Mux24~7_combout ),
	.datac(\storeregister[31][7]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~8 .lut_mask = 16'hE2CC;
defparam \Mux24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N23
dffeas \storeregister[22][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][7] .is_wysiwyg = "true";
defparam \storeregister[22][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N7
dffeas \storeregister[18][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][7] .is_wysiwyg = "true";
defparam \storeregister[18][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N6
cycloneive_lcell_comb \Mux24~2 (
// Equation(s):
// \Mux24~2_combout  = (temp_imemload_output_23 & ((\storeregister[22][7]~q ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\storeregister[18][7]~q  & !temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[22][7]~q ),
	.datac(\storeregister[18][7]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~2 .lut_mask = 16'hAAD8;
defparam \Mux24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N28
cycloneive_lcell_comb \storeregister[30][7]~feeder (
// Equation(s):
// \storeregister[30][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux24),
	.cin(gnd),
	.combout(\storeregister[30][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][7]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[30][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N29
dffeas \storeregister[30][7] (
	.clk(!CLK),
	.d(\storeregister[30][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][7] .is_wysiwyg = "true";
defparam \storeregister[30][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N30
cycloneive_lcell_comb \Mux24~3 (
// Equation(s):
// \Mux24~3_combout  = (temp_imemload_output_24 & ((\Mux24~2_combout  & ((\storeregister[30][7]~q ))) # (!\Mux24~2_combout  & (\storeregister[26][7]~q )))) # (!temp_imemload_output_24 & (((\Mux24~2_combout ))))

	.dataa(\storeregister[26][7]~q ),
	.datab(temp_imemload_output_24),
	.datac(\Mux24~2_combout ),
	.datad(\storeregister[30][7]~q ),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~3 .lut_mask = 16'hF838;
defparam \Mux24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N24
cycloneive_lcell_comb \storeregister[24][7]~feeder (
// Equation(s):
// \storeregister[24][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux24),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[24][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][7]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[24][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N25
dffeas \storeregister[24][7] (
	.clk(!CLK),
	.d(\storeregister[24][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][7] .is_wysiwyg = "true";
defparam \storeregister[24][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N31
dffeas \storeregister[28][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][7] .is_wysiwyg = "true";
defparam \storeregister[28][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N23
dffeas \storeregister[16][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][7] .is_wysiwyg = "true";
defparam \storeregister[16][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N6
cycloneive_lcell_comb \storeregister[20][7]~feeder (
// Equation(s):
// \storeregister[20][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux24),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[20][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][7]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[20][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N7
dffeas \storeregister[20][7] (
	.clk(!CLK),
	.d(\storeregister[20][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][7] .is_wysiwyg = "true";
defparam \storeregister[20][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N8
cycloneive_lcell_comb \Mux24~4 (
// Equation(s):
// \Mux24~4_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[20][7]~q ))) # (!temp_imemload_output_23 & (\storeregister[16][7]~q ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[16][7]~q ),
	.datac(temp_imemload_output_23),
	.datad(\storeregister[20][7]~q ),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~4 .lut_mask = 16'hF4A4;
defparam \Mux24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N12
cycloneive_lcell_comb \Mux24~5 (
// Equation(s):
// \Mux24~5_combout  = (temp_imemload_output_24 & ((\Mux24~4_combout  & ((\storeregister[28][7]~q ))) # (!\Mux24~4_combout  & (\storeregister[24][7]~q )))) # (!temp_imemload_output_24 & (((\Mux24~4_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[24][7]~q ),
	.datac(\storeregister[28][7]~q ),
	.datad(\Mux24~4_combout ),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~5 .lut_mask = 16'hF588;
defparam \Mux24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N16
cycloneive_lcell_comb \Mux24~6 (
// Equation(s):
// \Mux24~6_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\Mux24~3_combout )) # (!temp_imemload_output_22 & ((\Mux24~5_combout )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\Mux24~3_combout ),
	.datad(\Mux24~5_combout ),
	.cin(gnd),
	.combout(\Mux24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~6 .lut_mask = 16'hD9C8;
defparam \Mux24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N5
dffeas \storeregister[6][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][7] .is_wysiwyg = "true";
defparam \storeregister[6][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y41_N17
dffeas \storeregister[5][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][7] .is_wysiwyg = "true";
defparam \storeregister[5][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y41_N3
dffeas \storeregister[4][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][7] .is_wysiwyg = "true";
defparam \storeregister[4][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N16
cycloneive_lcell_comb \Mux24~10 (
// Equation(s):
// \Mux24~10_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[5][7]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[4][7]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[5][7]~q ),
	.datad(\storeregister[4][7]~q ),
	.cin(gnd),
	.combout(\Mux24~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~10 .lut_mask = 16'hB9A8;
defparam \Mux24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N12
cycloneive_lcell_comb \storeregister[7][7]~feeder (
// Equation(s):
// \storeregister[7][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux24),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[7][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[7][7]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[7][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N13
dffeas \storeregister[7][7] (
	.clk(!CLK),
	.d(\storeregister[7][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][7] .is_wysiwyg = "true";
defparam \storeregister[7][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N14
cycloneive_lcell_comb \Mux24~11 (
// Equation(s):
// \Mux24~11_combout  = (temp_imemload_output_22 & ((\Mux24~10_combout  & ((\storeregister[7][7]~q ))) # (!\Mux24~10_combout  & (\storeregister[6][7]~q )))) # (!temp_imemload_output_22 & (((\Mux24~10_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[6][7]~q ),
	.datac(\Mux24~10_combout ),
	.datad(\storeregister[7][7]~q ),
	.cin(gnd),
	.combout(\Mux24~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~11 .lut_mask = 16'hF858;
defparam \Mux24~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N12
cycloneive_lcell_comb \storeregister[14][7]~feeder (
// Equation(s):
// \storeregister[14][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux24),
	.cin(gnd),
	.combout(\storeregister[14][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][7]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N13
dffeas \storeregister[14][7] (
	.clk(!CLK),
	.d(\storeregister[14][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][7] .is_wysiwyg = "true";
defparam \storeregister[14][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N5
dffeas \storeregister[15][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][7] .is_wysiwyg = "true";
defparam \storeregister[15][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N27
dffeas \storeregister[13][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][7] .is_wysiwyg = "true";
defparam \storeregister[13][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N1
dffeas \storeregister[12][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][7] .is_wysiwyg = "true";
defparam \storeregister[12][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N26
cycloneive_lcell_comb \Mux24~17 (
// Equation(s):
// \Mux24~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][7]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[12][7]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[13][7]~q ),
	.datad(\storeregister[12][7]~q ),
	.cin(gnd),
	.combout(\Mux24~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~17 .lut_mask = 16'hB9A8;
defparam \Mux24~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N26
cycloneive_lcell_comb \Mux24~18 (
// Equation(s):
// \Mux24~18_combout  = (temp_imemload_output_22 & ((\Mux24~17_combout  & ((\storeregister[15][7]~q ))) # (!\Mux24~17_combout  & (\storeregister[14][7]~q )))) # (!temp_imemload_output_22 & (((\Mux24~17_combout ))))

	.dataa(\storeregister[14][7]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[15][7]~q ),
	.datad(\Mux24~17_combout ),
	.cin(gnd),
	.combout(\Mux24~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~18 .lut_mask = 16'hF388;
defparam \Mux24~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N19
dffeas \storeregister[8][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][7] .is_wysiwyg = "true";
defparam \storeregister[8][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N21
dffeas \storeregister[10][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][7] .is_wysiwyg = "true";
defparam \storeregister[10][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N18
cycloneive_lcell_comb \Mux24~12 (
// Equation(s):
// \Mux24~12_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\storeregister[10][7]~q )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & (\storeregister[8][7]~q )))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[8][7]~q ),
	.datad(\storeregister[10][7]~q ),
	.cin(gnd),
	.combout(\Mux24~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~12 .lut_mask = 16'hBA98;
defparam \Mux24~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N24
cycloneive_lcell_comb \storeregister[9][7]~feeder (
// Equation(s):
// \storeregister[9][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux24),
	.cin(gnd),
	.combout(\storeregister[9][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[9][7]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[9][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N25
dffeas \storeregister[9][7] (
	.clk(!CLK),
	.d(\storeregister[9][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][7] .is_wysiwyg = "true";
defparam \storeregister[9][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N16
cycloneive_lcell_comb \Mux24~13 (
// Equation(s):
// \Mux24~13_combout  = (temp_imemload_output_21 & ((\Mux24~12_combout  & (\storeregister[11][7]~q )) # (!\Mux24~12_combout  & ((\storeregister[9][7]~q ))))) # (!temp_imemload_output_21 & (((\Mux24~12_combout ))))

	.dataa(\storeregister[11][7]~q ),
	.datab(temp_imemload_output_21),
	.datac(\Mux24~12_combout ),
	.datad(\storeregister[9][7]~q ),
	.cin(gnd),
	.combout(\Mux24~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~13 .lut_mask = 16'hBCB0;
defparam \Mux24~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N5
dffeas \storeregister[3][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][7] .is_wysiwyg = "true";
defparam \storeregister[3][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N19
dffeas \storeregister[1][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][7] .is_wysiwyg = "true";
defparam \storeregister[1][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N18
cycloneive_lcell_comb \Mux24~14 (
// Equation(s):
// \Mux24~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[3][7]~q )) # (!temp_imemload_output_22 & ((\storeregister[1][7]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[3][7]~q ),
	.datac(\storeregister[1][7]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux24~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~14 .lut_mask = 16'h88A0;
defparam \Mux24~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N27
dffeas \storeregister[2][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][7] .is_wysiwyg = "true";
defparam \storeregister[2][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N20
cycloneive_lcell_comb \Mux24~15 (
// Equation(s):
// \Mux24~15_combout  = (\Mux24~14_combout ) # ((!temp_imemload_output_21 & (\storeregister[2][7]~q  & temp_imemload_output_22)))

	.dataa(temp_imemload_output_21),
	.datab(\Mux24~14_combout ),
	.datac(\storeregister[2][7]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux24~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~15 .lut_mask = 16'hDCCC;
defparam \Mux24~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N12
cycloneive_lcell_comb \Mux24~16 (
// Equation(s):
// \Mux24~16_combout  = (temp_imemload_output_24 & ((\Mux24~13_combout ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((!temp_imemload_output_23 & \Mux24~15_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\Mux24~13_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux24~15_combout ),
	.cin(gnd),
	.combout(\Mux24~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~16 .lut_mask = 16'hADA8;
defparam \Mux24~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N4
cycloneive_lcell_comb \storeregister[28][6]~feeder (
// Equation(s):
// \storeregister[28][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux25),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[28][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][6]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[28][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N5
dffeas \storeregister[28][6] (
	.clk(!CLK),
	.d(\storeregister[28][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][6] .is_wysiwyg = "true";
defparam \storeregister[28][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N8
cycloneive_lcell_comb \storeregister[16][6]~feeder (
// Equation(s):
// \storeregister[16][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux25),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[16][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[16][6]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[16][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N9
dffeas \storeregister[16][6] (
	.clk(!CLK),
	.d(\storeregister[16][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][6] .is_wysiwyg = "true";
defparam \storeregister[16][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N16
cycloneive_lcell_comb \storeregister[24][6]~feeder (
// Equation(s):
// \storeregister[24][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux25),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[24][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][6]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[24][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N17
dffeas \storeregister[24][6] (
	.clk(!CLK),
	.d(\storeregister[24][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][6] .is_wysiwyg = "true";
defparam \storeregister[24][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N6
cycloneive_lcell_comb \Mux25~4 (
// Equation(s):
// \Mux25~4_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[24][6]~q ))) # (!temp_imemload_output_24 & (\storeregister[16][6]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][6]~q ),
	.datad(\storeregister[24][6]~q ),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~4 .lut_mask = 16'hDC98;
defparam \Mux25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N2
cycloneive_lcell_comb \storeregister[20][6]~feeder (
// Equation(s):
// \storeregister[20][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux25),
	.cin(gnd),
	.combout(\storeregister[20][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][6]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[20][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N3
dffeas \storeregister[20][6] (
	.clk(!CLK),
	.d(\storeregister[20][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][6] .is_wysiwyg = "true";
defparam \storeregister[20][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N4
cycloneive_lcell_comb \Mux25~5 (
// Equation(s):
// \Mux25~5_combout  = (temp_imemload_output_23 & ((\Mux25~4_combout  & (\storeregister[28][6]~q )) # (!\Mux25~4_combout  & ((\storeregister[20][6]~q ))))) # (!temp_imemload_output_23 & (((\Mux25~4_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[28][6]~q ),
	.datac(\Mux25~4_combout ),
	.datad(\storeregister[20][6]~q ),
	.cin(gnd),
	.combout(\Mux25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~5 .lut_mask = 16'hDAD0;
defparam \Mux25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N29
dffeas \storeregister[22][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][6] .is_wysiwyg = "true";
defparam \storeregister[22][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N15
dffeas \storeregister[30][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][6] .is_wysiwyg = "true";
defparam \storeregister[30][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N1
dffeas \storeregister[26][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][6] .is_wysiwyg = "true";
defparam \storeregister[26][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N11
dffeas \storeregister[18][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][6] .is_wysiwyg = "true";
defparam \storeregister[18][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N10
cycloneive_lcell_comb \Mux25~2 (
// Equation(s):
// \Mux25~2_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[26][6]~q )) # (!temp_imemload_output_24 & ((\storeregister[18][6]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[26][6]~q ),
	.datac(\storeregister[18][6]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~2 .lut_mask = 16'hEE50;
defparam \Mux25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N14
cycloneive_lcell_comb \Mux25~3 (
// Equation(s):
// \Mux25~3_combout  = (temp_imemload_output_23 & ((\Mux25~2_combout  & ((\storeregister[30][6]~q ))) # (!\Mux25~2_combout  & (\storeregister[22][6]~q )))) # (!temp_imemload_output_23 & (((\Mux25~2_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[22][6]~q ),
	.datac(\storeregister[30][6]~q ),
	.datad(\Mux25~2_combout ),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~3 .lut_mask = 16'hF588;
defparam \Mux25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N6
cycloneive_lcell_comb \Mux25~6 (
// Equation(s):
// \Mux25~6_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\Mux25~3_combout )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & (\Mux25~5_combout )))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\Mux25~5_combout ),
	.datad(\Mux25~3_combout ),
	.cin(gnd),
	.combout(\Mux25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~6 .lut_mask = 16'hBA98;
defparam \Mux25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N4
cycloneive_lcell_comb \storeregister[23][6]~feeder (
// Equation(s):
// \storeregister[23][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux25),
	.cin(gnd),
	.combout(\storeregister[23][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][6]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[23][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N5
dffeas \storeregister[23][6] (
	.clk(!CLK),
	.d(\storeregister[23][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][6] .is_wysiwyg = "true";
defparam \storeregister[23][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N18
cycloneive_lcell_comb \storeregister[19][6]~feeder (
// Equation(s):
// \storeregister[19][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux25),
	.cin(gnd),
	.combout(\storeregister[19][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[19][6]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[19][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N19
dffeas \storeregister[19][6] (
	.clk(!CLK),
	.d(\storeregister[19][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][6] .is_wysiwyg = "true";
defparam \storeregister[19][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N12
cycloneive_lcell_comb \Mux25~7 (
// Equation(s):
// \Mux25~7_combout  = (temp_imemload_output_23 & ((\storeregister[23][6]~q ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((!temp_imemload_output_24 & \storeregister[19][6]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[23][6]~q ),
	.datac(temp_imemload_output_24),
	.datad(\storeregister[19][6]~q ),
	.cin(gnd),
	.combout(\Mux25~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~7 .lut_mask = 16'hADA8;
defparam \Mux25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N12
cycloneive_lcell_comb \storeregister[27][6]~feeder (
// Equation(s):
// \storeregister[27][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux25),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][6]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N13
dffeas \storeregister[27][6] (
	.clk(!CLK),
	.d(\storeregister[27][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][6] .is_wysiwyg = "true";
defparam \storeregister[27][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N6
cycloneive_lcell_comb \storeregister[31][6]~feeder (
// Equation(s):
// \storeregister[31][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux25),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[31][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][6]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[31][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N7
dffeas \storeregister[31][6] (
	.clk(!CLK),
	.d(\storeregister[31][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][6] .is_wysiwyg = "true";
defparam \storeregister[31][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N18
cycloneive_lcell_comb \Mux25~8 (
// Equation(s):
// \Mux25~8_combout  = (\Mux25~7_combout  & (((\storeregister[31][6]~q ) # (!temp_imemload_output_24)))) # (!\Mux25~7_combout  & (\storeregister[27][6]~q  & (temp_imemload_output_24)))

	.dataa(\Mux25~7_combout ),
	.datab(\storeregister[27][6]~q ),
	.datac(temp_imemload_output_24),
	.datad(\storeregister[31][6]~q ),
	.cin(gnd),
	.combout(\Mux25~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~8 .lut_mask = 16'hEA4A;
defparam \Mux25~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N25
dffeas \storeregister[21][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][6] .is_wysiwyg = "true";
defparam \storeregister[21][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N24
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (temp_imemload_output_23 & (((\storeregister[21][6]~q ) # (temp_imemload_output_24)))) # (!temp_imemload_output_23 & (\storeregister[17][6]~q  & ((!temp_imemload_output_24))))

	.dataa(\storeregister[17][6]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[21][6]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hCCE2;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N29
dffeas \storeregister[25][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][6] .is_wysiwyg = "true";
defparam \storeregister[25][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N28
cycloneive_lcell_comb \storeregister[29][6]~feeder (
// Equation(s):
// \storeregister[29][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux25),
	.cin(gnd),
	.combout(\storeregister[29][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][6]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[29][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y42_N29
dffeas \storeregister[29][6] (
	.clk(!CLK),
	.d(\storeregister[29][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][6] .is_wysiwyg = "true";
defparam \storeregister[29][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N28
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\Mux25~0_combout  & (((\storeregister[29][6]~q )) # (!temp_imemload_output_24))) # (!\Mux25~0_combout  & (temp_imemload_output_24 & (\storeregister[25][6]~q )))

	.dataa(\Mux25~0_combout ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[25][6]~q ),
	.datad(\storeregister[29][6]~q ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hEA62;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N27
dffeas \storeregister[11][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][6] .is_wysiwyg = "true";
defparam \storeregister[11][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N21
dffeas \storeregister[10][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][6] .is_wysiwyg = "true";
defparam \storeregister[10][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N29
dffeas \storeregister[8][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][6] .is_wysiwyg = "true";
defparam \storeregister[8][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N20
cycloneive_lcell_comb \Mux25~10 (
// Equation(s):
// \Mux25~10_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[10][6]~q )) # (!temp_imemload_output_22 & ((\storeregister[8][6]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][6]~q ),
	.datad(\storeregister[8][6]~q ),
	.cin(gnd),
	.combout(\Mux25~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~10 .lut_mask = 16'hD9C8;
defparam \Mux25~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N3
dffeas \storeregister[9][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][6] .is_wysiwyg = "true";
defparam \storeregister[9][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N2
cycloneive_lcell_comb \Mux25~11 (
// Equation(s):
// \Mux25~11_combout  = (\Mux25~10_combout  & ((\storeregister[11][6]~q ) # ((!temp_imemload_output_21)))) # (!\Mux25~10_combout  & (((\storeregister[9][6]~q  & temp_imemload_output_21))))

	.dataa(\storeregister[11][6]~q ),
	.datab(\Mux25~10_combout ),
	.datac(\storeregister[9][6]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux25~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~11 .lut_mask = 16'hB8CC;
defparam \Mux25~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N3
dffeas \storeregister[7][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][6] .is_wysiwyg = "true";
defparam \storeregister[7][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N25
dffeas \storeregister[6][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][6] .is_wysiwyg = "true";
defparam \storeregister[6][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N2
cycloneive_lcell_comb \Mux25~13 (
// Equation(s):
// \Mux25~13_combout  = (\Mux25~12_combout  & (((\storeregister[7][6]~q )) # (!temp_imemload_output_22))) # (!\Mux25~12_combout  & (temp_imemload_output_22 & ((\storeregister[6][6]~q ))))

	.dataa(\Mux25~12_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[7][6]~q ),
	.datad(\storeregister[6][6]~q ),
	.cin(gnd),
	.combout(\Mux25~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~13 .lut_mask = 16'hE6A2;
defparam \Mux25~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N25
dffeas \storeregister[3][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][6] .is_wysiwyg = "true";
defparam \storeregister[3][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N11
dffeas \storeregister[1][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][6] .is_wysiwyg = "true";
defparam \storeregister[1][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N10
cycloneive_lcell_comb \Mux25~14 (
// Equation(s):
// \Mux25~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[3][6]~q )) # (!temp_imemload_output_22 & ((\storeregister[1][6]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[3][6]~q ),
	.datac(\storeregister[1][6]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux25~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~14 .lut_mask = 16'h88A0;
defparam \Mux25~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N8
cycloneive_lcell_comb \storeregister[2][6]~feeder (
// Equation(s):
// \storeregister[2][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux25),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[2][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[2][6]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[2][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N9
dffeas \storeregister[2][6] (
	.clk(!CLK),
	.d(\storeregister[2][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][6] .is_wysiwyg = "true";
defparam \storeregister[2][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N20
cycloneive_lcell_comb \Mux25~15 (
// Equation(s):
// \Mux25~15_combout  = (\Mux25~14_combout ) # ((temp_imemload_output_22 & (!temp_imemload_output_21 & \storeregister[2][6]~q )))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\Mux25~14_combout ),
	.datad(\storeregister[2][6]~q ),
	.cin(gnd),
	.combout(\Mux25~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~15 .lut_mask = 16'hF2F0;
defparam \Mux25~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N6
cycloneive_lcell_comb \Mux25~16 (
// Equation(s):
// \Mux25~16_combout  = (temp_imemload_output_23 & ((\Mux25~13_combout ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\Mux25~15_combout  & !temp_imemload_output_24))))

	.dataa(\Mux25~13_combout ),
	.datab(\Mux25~15_combout ),
	.datac(temp_imemload_output_23),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux25~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~16 .lut_mask = 16'hF0AC;
defparam \Mux25~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N30
cycloneive_lcell_comb \storeregister[15][6]~feeder (
// Equation(s):
// \storeregister[15][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux25),
	.cin(gnd),
	.combout(\storeregister[15][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][6]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y44_N31
dffeas \storeregister[15][6] (
	.clk(!CLK),
	.d(\storeregister[15][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][6] .is_wysiwyg = "true";
defparam \storeregister[15][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N3
dffeas \storeregister[13][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][6] .is_wysiwyg = "true";
defparam \storeregister[13][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N17
dffeas \storeregister[12][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][6] .is_wysiwyg = "true";
defparam \storeregister[12][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N2
cycloneive_lcell_comb \Mux25~17 (
// Equation(s):
// \Mux25~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][6]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[12][6]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[13][6]~q ),
	.datad(\storeregister[12][6]~q ),
	.cin(gnd),
	.combout(\Mux25~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~17 .lut_mask = 16'hB9A8;
defparam \Mux25~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N8
cycloneive_lcell_comb \storeregister[14][6]~feeder (
// Equation(s):
// \storeregister[14][6]~feeder_combout  = Mux25

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux25),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[14][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][6]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[14][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N9
dffeas \storeregister[14][6] (
	.clk(!CLK),
	.d(\storeregister[14][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][6] .is_wysiwyg = "true";
defparam \storeregister[14][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N18
cycloneive_lcell_comb \Mux25~18 (
// Equation(s):
// \Mux25~18_combout  = (\Mux25~17_combout  & ((\storeregister[15][6]~q ) # ((!temp_imemload_output_22)))) # (!\Mux25~17_combout  & (((\storeregister[14][6]~q  & temp_imemload_output_22))))

	.dataa(\storeregister[15][6]~q ),
	.datab(\Mux25~17_combout ),
	.datac(\storeregister[14][6]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux25~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~18 .lut_mask = 16'hB8CC;
defparam \Mux25~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N30
cycloneive_lcell_comb \storeregister[18][5]~feeder (
// Equation(s):
// \storeregister[18][5]~feeder_combout  = Mux26

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux26),
	.cin(gnd),
	.combout(\storeregister[18][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[18][5]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[18][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N31
dffeas \storeregister[18][5] (
	.clk(!CLK),
	.d(\storeregister[18][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][5] .is_wysiwyg = "true";
defparam \storeregister[18][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N8
cycloneive_lcell_comb \Mux26~2 (
// Equation(s):
// \Mux26~2_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[22][5]~q )) # (!temp_imemload_output_23 & ((\storeregister[18][5]~q )))))

	.dataa(\storeregister[22][5]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[18][5]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~2 .lut_mask = 16'hEE30;
defparam \Mux26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N0
cycloneive_lcell_comb \storeregister[26][5]~feeder (
// Equation(s):
// \storeregister[26][5]~feeder_combout  = Mux26

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux26),
	.cin(gnd),
	.combout(\storeregister[26][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[26][5]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[26][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N1
dffeas \storeregister[26][5] (
	.clk(!CLK),
	.d(\storeregister[26][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][5] .is_wysiwyg = "true";
defparam \storeregister[26][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N6
cycloneive_lcell_comb \Mux26~3 (
// Equation(s):
// \Mux26~3_combout  = (temp_imemload_output_24 & ((\Mux26~2_combout  & (\storeregister[30][5]~q )) # (!\Mux26~2_combout  & ((\storeregister[26][5]~q ))))) # (!temp_imemload_output_24 & (((\Mux26~2_combout ))))

	.dataa(\storeregister[30][5]~q ),
	.datab(temp_imemload_output_24),
	.datac(\Mux26~2_combout ),
	.datad(\storeregister[26][5]~q ),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~3 .lut_mask = 16'hBCB0;
defparam \Mux26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N29
dffeas \storeregister[28][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][5] .is_wysiwyg = "true";
defparam \storeregister[28][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N24
cycloneive_lcell_comb \storeregister[20][5]~feeder (
// Equation(s):
// \storeregister[20][5]~feeder_combout  = Mux26

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux26),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[20][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][5]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[20][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N25
dffeas \storeregister[20][5] (
	.clk(!CLK),
	.d(\storeregister[20][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][5] .is_wysiwyg = "true";
defparam \storeregister[20][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N6
cycloneive_lcell_comb \Mux26~4 (
// Equation(s):
// \Mux26~4_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24) # (\storeregister[20][5]~q )))) # (!temp_imemload_output_23 & (\storeregister[16][5]~q  & (!temp_imemload_output_24)))

	.dataa(\storeregister[16][5]~q ),
	.datab(temp_imemload_output_23),
	.datac(temp_imemload_output_24),
	.datad(\storeregister[20][5]~q ),
	.cin(gnd),
	.combout(\Mux26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~4 .lut_mask = 16'hCEC2;
defparam \Mux26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N28
cycloneive_lcell_comb \Mux26~5 (
// Equation(s):
// \Mux26~5_combout  = (temp_imemload_output_24 & ((\Mux26~4_combout  & ((\storeregister[28][5]~q ))) # (!\Mux26~4_combout  & (\storeregister[24][5]~q )))) # (!temp_imemload_output_24 & (((\Mux26~4_combout ))))

	.dataa(\storeregister[24][5]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[28][5]~q ),
	.datad(\Mux26~4_combout ),
	.cin(gnd),
	.combout(\Mux26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~5 .lut_mask = 16'hF388;
defparam \Mux26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N16
cycloneive_lcell_comb \Mux26~6 (
// Equation(s):
// \Mux26~6_combout  = (temp_imemload_output_22 & ((\Mux26~3_combout ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((\Mux26~5_combout  & !temp_imemload_output_21))))

	.dataa(\Mux26~3_combout ),
	.datab(\Mux26~5_combout ),
	.datac(temp_imemload_output_22),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~6 .lut_mask = 16'hF0AC;
defparam \Mux26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N15
dffeas \storeregister[31][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][5] .is_wysiwyg = "true";
defparam \storeregister[31][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N25
dffeas \storeregister[23][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][5] .is_wysiwyg = "true";
defparam \storeregister[23][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N31
dffeas \storeregister[19][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][5] .is_wysiwyg = "true";
defparam \storeregister[19][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N29
dffeas \storeregister[27][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][5] .is_wysiwyg = "true";
defparam \storeregister[27][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N28
cycloneive_lcell_comb \Mux26~7 (
// Equation(s):
// \Mux26~7_combout  = (temp_imemload_output_24 & (((\storeregister[27][5]~q ) # (temp_imemload_output_23)))) # (!temp_imemload_output_24 & (\storeregister[19][5]~q  & ((!temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[19][5]~q ),
	.datac(\storeregister[27][5]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux26~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~7 .lut_mask = 16'hAAE4;
defparam \Mux26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N24
cycloneive_lcell_comb \Mux26~8 (
// Equation(s):
// \Mux26~8_combout  = (temp_imemload_output_23 & ((\Mux26~7_combout  & (\storeregister[31][5]~q )) # (!\Mux26~7_combout  & ((\storeregister[23][5]~q ))))) # (!temp_imemload_output_23 & (((\Mux26~7_combout ))))

	.dataa(\storeregister[31][5]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[23][5]~q ),
	.datad(\Mux26~7_combout ),
	.cin(gnd),
	.combout(\Mux26~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~8 .lut_mask = 16'hBBC0;
defparam \Mux26~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N20
cycloneive_lcell_comb \storeregister[17][5]~feeder (
// Equation(s):
// \storeregister[17][5]~feeder_combout  = Mux26

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux26),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[17][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[17][5]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[17][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N21
dffeas \storeregister[17][5] (
	.clk(!CLK),
	.d(\storeregister[17][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][5] .is_wysiwyg = "true";
defparam \storeregister[17][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N4
cycloneive_lcell_comb \storeregister[25][5]~feeder (
// Equation(s):
// \storeregister[25][5]~feeder_combout  = Mux26

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux26),
	.cin(gnd),
	.combout(\storeregister[25][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[25][5]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[25][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N5
dffeas \storeregister[25][5] (
	.clk(!CLK),
	.d(\storeregister[25][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][5] .is_wysiwyg = "true";
defparam \storeregister[25][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N30
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (temp_imemload_output_24 & (((\storeregister[25][5]~q ) # (temp_imemload_output_23)))) # (!temp_imemload_output_24 & (\storeregister[17][5]~q  & ((!temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[17][5]~q ),
	.datac(\storeregister[25][5]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hAAE4;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N20
cycloneive_lcell_comb \storeregister[21][5]~feeder (
// Equation(s):
// \storeregister[21][5]~feeder_combout  = Mux26

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux26),
	.cin(gnd),
	.combout(\storeregister[21][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][5]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[21][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N21
dffeas \storeregister[21][5] (
	.clk(!CLK),
	.d(\storeregister[21][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][5] .is_wysiwyg = "true";
defparam \storeregister[21][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N30
cycloneive_lcell_comb \storeregister[29][5]~feeder (
// Equation(s):
// \storeregister[29][5]~feeder_combout  = Mux26

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux26),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[29][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][5]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[29][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N31
dffeas \storeregister[29][5] (
	.clk(!CLK),
	.d(\storeregister[29][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][5] .is_wysiwyg = "true";
defparam \storeregister[29][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N10
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (\Mux26~0_combout  & (((\storeregister[29][5]~q )) # (!temp_imemload_output_23))) # (!\Mux26~0_combout  & (temp_imemload_output_23 & (\storeregister[21][5]~q )))

	.dataa(\Mux26~0_combout ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[21][5]~q ),
	.datad(\storeregister[29][5]~q ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hEA62;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N7
dffeas \storeregister[11][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][5] .is_wysiwyg = "true";
defparam \storeregister[11][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N29
dffeas \storeregister[9][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][5] .is_wysiwyg = "true";
defparam \storeregister[9][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N6
cycloneive_lcell_comb \Mux26~13 (
// Equation(s):
// \Mux26~13_combout  = (\Mux26~12_combout  & (((\storeregister[11][5]~q )) # (!temp_imemload_output_21))) # (!\Mux26~12_combout  & (temp_imemload_output_21 & ((\storeregister[9][5]~q ))))

	.dataa(\Mux26~12_combout ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[11][5]~q ),
	.datad(\storeregister[9][5]~q ),
	.cin(gnd),
	.combout(\Mux26~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~13 .lut_mask = 16'hE6A2;
defparam \Mux26~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N15
dffeas \storeregister[2][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][5] .is_wysiwyg = "true";
defparam \storeregister[2][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N15
dffeas \storeregister[1][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][5] .is_wysiwyg = "true";
defparam \storeregister[1][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N29
dffeas \storeregister[3][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][5] .is_wysiwyg = "true";
defparam \storeregister[3][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N14
cycloneive_lcell_comb \Mux26~14 (
// Equation(s):
// \Mux26~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][5]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][5]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[1][5]~q ),
	.datad(\storeregister[3][5]~q ),
	.cin(gnd),
	.combout(\Mux26~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~14 .lut_mask = 16'hA820;
defparam \Mux26~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N18
cycloneive_lcell_comb \Mux26~15 (
// Equation(s):
// \Mux26~15_combout  = (\Mux26~14_combout ) # ((!temp_imemload_output_21 & (\storeregister[2][5]~q  & temp_imemload_output_22)))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[2][5]~q ),
	.datac(temp_imemload_output_22),
	.datad(\Mux26~14_combout ),
	.cin(gnd),
	.combout(\Mux26~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~15 .lut_mask = 16'hFF40;
defparam \Mux26~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N4
cycloneive_lcell_comb \Mux26~16 (
// Equation(s):
// \Mux26~16_combout  = (temp_imemload_output_24 & ((temp_imemload_output_23) # ((\Mux26~13_combout )))) # (!temp_imemload_output_24 & (!temp_imemload_output_23 & ((\Mux26~15_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\Mux26~13_combout ),
	.datad(\Mux26~15_combout ),
	.cin(gnd),
	.combout(\Mux26~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~16 .lut_mask = 16'hB9A8;
defparam \Mux26~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N10
cycloneive_lcell_comb \storeregister[14][5]~feeder (
// Equation(s):
// \storeregister[14][5]~feeder_combout  = Mux26

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux26),
	.cin(gnd),
	.combout(\storeregister[14][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][5]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N11
dffeas \storeregister[14][5] (
	.clk(!CLK),
	.d(\storeregister[14][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][5] .is_wysiwyg = "true";
defparam \storeregister[14][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N8
cycloneive_lcell_comb \storeregister[15][5]~feeder (
// Equation(s):
// \storeregister[15][5]~feeder_combout  = Mux26

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux26),
	.cin(gnd),
	.combout(\storeregister[15][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][5]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N9
dffeas \storeregister[15][5] (
	.clk(!CLK),
	.d(\storeregister[15][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][5] .is_wysiwyg = "true";
defparam \storeregister[15][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N31
dffeas \storeregister[13][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][5] .is_wysiwyg = "true";
defparam \storeregister[13][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N13
dffeas \storeregister[12][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][5] .is_wysiwyg = "true";
defparam \storeregister[12][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N30
cycloneive_lcell_comb \Mux26~17 (
// Equation(s):
// \Mux26~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][5]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[12][5]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[13][5]~q ),
	.datad(\storeregister[12][5]~q ),
	.cin(gnd),
	.combout(\Mux26~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~17 .lut_mask = 16'hB9A8;
defparam \Mux26~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N30
cycloneive_lcell_comb \Mux26~18 (
// Equation(s):
// \Mux26~18_combout  = (\Mux26~17_combout  & (((\storeregister[15][5]~q ) # (!temp_imemload_output_22)))) # (!\Mux26~17_combout  & (\storeregister[14][5]~q  & ((temp_imemload_output_22))))

	.dataa(\storeregister[14][5]~q ),
	.datab(\storeregister[15][5]~q ),
	.datac(\Mux26~17_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux26~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~18 .lut_mask = 16'hCAF0;
defparam \Mux26~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y41_N13
dffeas \storeregister[5][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][5] .is_wysiwyg = "true";
defparam \storeregister[5][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y41_N27
dffeas \storeregister[4][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][5] .is_wysiwyg = "true";
defparam \storeregister[4][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N12
cycloneive_lcell_comb \Mux26~10 (
// Equation(s):
// \Mux26~10_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[5][5]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[4][5]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[5][5]~q ),
	.datad(\storeregister[4][5]~q ),
	.cin(gnd),
	.combout(\Mux26~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~10 .lut_mask = 16'hB9A8;
defparam \Mux26~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N17
dffeas \storeregister[7][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][5] .is_wysiwyg = "true";
defparam \storeregister[7][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N7
dffeas \storeregister[6][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][5] .is_wysiwyg = "true";
defparam \storeregister[6][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N6
cycloneive_lcell_comb \Mux26~11 (
// Equation(s):
// \Mux26~11_combout  = (\Mux26~10_combout  & ((\storeregister[7][5]~q ) # ((!temp_imemload_output_22)))) # (!\Mux26~10_combout  & (((\storeregister[6][5]~q  & temp_imemload_output_22))))

	.dataa(\Mux26~10_combout ),
	.datab(\storeregister[7][5]~q ),
	.datac(\storeregister[6][5]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux26~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~11 .lut_mask = 16'hD8AA;
defparam \Mux26~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N24
cycloneive_lcell_comb \storeregister[24][3]~feeder (
// Equation(s):
// \storeregister[24][3]~feeder_combout  = Mux28

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux28),
	.cin(gnd),
	.combout(\storeregister[24][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][3]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[24][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N25
dffeas \storeregister[24][3] (
	.clk(!CLK),
	.d(\storeregister[24][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][3] .is_wysiwyg = "true";
defparam \storeregister[24][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N18
cycloneive_lcell_comb \Mux60~4 (
// Equation(s):
// \Mux60~4_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\storeregister[24][3]~q )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & (\storeregister[16][3]~q )))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[16][3]~q ),
	.datad(\storeregister[24][3]~q ),
	.cin(gnd),
	.combout(\Mux60~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~4 .lut_mask = 16'hBA98;
defparam \Mux60~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N28
cycloneive_lcell_comb \Mux60~5 (
// Equation(s):
// \Mux60~5_combout  = (temp_imemload_output_18 & ((\Mux60~4_combout  & (\storeregister[28][3]~q )) # (!\Mux60~4_combout  & ((\storeregister[20][3]~q ))))) # (!temp_imemload_output_18 & (\Mux60~4_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux60~4_combout ),
	.datac(\storeregister[28][3]~q ),
	.datad(\storeregister[20][3]~q ),
	.cin(gnd),
	.combout(\Mux60~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~5 .lut_mask = 16'hE6C4;
defparam \Mux60~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N16
cycloneive_lcell_comb \Mux60~2 (
// Equation(s):
// \Mux60~2_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\storeregister[26][3]~q )) # (!temp_imemload_output_19 & ((\storeregister[18][3]~q )))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[26][3]~q ),
	.datad(\storeregister[18][3]~q ),
	.cin(gnd),
	.combout(\Mux60~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~2 .lut_mask = 16'hD9C8;
defparam \Mux60~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N0
cycloneive_lcell_comb \Mux60~3 (
// Equation(s):
// \Mux60~3_combout  = (\Mux60~2_combout  & ((\storeregister[30][3]~q ) # ((!temp_imemload_output_18)))) # (!\Mux60~2_combout  & (((\storeregister[22][3]~q  & temp_imemload_output_18))))

	.dataa(\storeregister[30][3]~q ),
	.datab(\storeregister[22][3]~q ),
	.datac(\Mux60~2_combout ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux60~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~3 .lut_mask = 16'hACF0;
defparam \Mux60~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N20
cycloneive_lcell_comb \Mux60~6 (
// Equation(s):
// \Mux60~6_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16) # (\Mux60~3_combout )))) # (!temp_imemload_output_17 & (\Mux60~5_combout  & (!temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux60~5_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux60~3_combout ),
	.cin(gnd),
	.combout(\Mux60~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~6 .lut_mask = 16'hAEA4;
defparam \Mux60~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N28
cycloneive_lcell_comb \Mux60~0 (
// Equation(s):
// \Mux60~0_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[21][3]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[17][3]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[21][3]~q ),
	.datad(\storeregister[17][3]~q ),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~0 .lut_mask = 16'hB9A8;
defparam \Mux60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N18
cycloneive_lcell_comb \Mux60~1 (
// Equation(s):
// \Mux60~1_combout  = (\Mux60~0_combout  & (((\storeregister[29][3]~q ) # (!temp_imemload_output_19)))) # (!\Mux60~0_combout  & (\storeregister[25][3]~q  & (temp_imemload_output_19)))

	.dataa(\Mux60~0_combout ),
	.datab(\storeregister[25][3]~q ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[29][3]~q ),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~1 .lut_mask = 16'hEA4A;
defparam \Mux60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N3
dffeas \storeregister[19][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][3] .is_wysiwyg = "true";
defparam \storeregister[19][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N2
cycloneive_lcell_comb \Mux60~7 (
// Equation(s):
// \Mux60~7_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\storeregister[23][3]~q )) # (!temp_imemload_output_18 & ((\storeregister[19][3]~q )))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[23][3]~q ),
	.datac(\storeregister[19][3]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux60~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~7 .lut_mask = 16'hEE50;
defparam \Mux60~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N22
cycloneive_lcell_comb \Mux60~8 (
// Equation(s):
// \Mux60~8_combout  = (\Mux60~7_combout  & (((\storeregister[31][3]~q )) # (!temp_imemload_output_19))) # (!\Mux60~7_combout  & (temp_imemload_output_19 & (\storeregister[27][3]~q )))

	.dataa(\Mux60~7_combout ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[27][3]~q ),
	.datad(\storeregister[31][3]~q ),
	.cin(gnd),
	.combout(\Mux60~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~8 .lut_mask = 16'hEA62;
defparam \Mux60~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N10
cycloneive_lcell_comb \Mux60~12 (
// Equation(s):
// \Mux60~12_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[5][3]~q )) # (!temp_imemload_output_16 & ((\storeregister[4][3]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[5][3]~q ),
	.datac(\storeregister[4][3]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux60~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~12 .lut_mask = 16'hEE50;
defparam \Mux60~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N16
cycloneive_lcell_comb \Mux60~13 (
// Equation(s):
// \Mux60~13_combout  = (\Mux60~12_combout  & ((\storeregister[7][3]~q ) # ((!temp_imemload_output_17)))) # (!\Mux60~12_combout  & (((temp_imemload_output_17 & \storeregister[6][3]~q ))))

	.dataa(\storeregister[7][3]~q ),
	.datab(\Mux60~12_combout ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[6][3]~q ),
	.cin(gnd),
	.combout(\Mux60~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~13 .lut_mask = 16'hBC8C;
defparam \Mux60~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N15
dffeas \storeregister[1][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][3] .is_wysiwyg = "true";
defparam \storeregister[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N1
dffeas \storeregister[3][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][3] .is_wysiwyg = "true";
defparam \storeregister[3][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N0
cycloneive_lcell_comb \Mux60~14 (
// Equation(s):
// \Mux60~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[3][3]~q ))) # (!temp_imemload_output_17 & (\storeregister[1][3]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[1][3]~q ),
	.datac(\storeregister[3][3]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux60~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~14 .lut_mask = 16'hA088;
defparam \Mux60~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N30
cycloneive_lcell_comb \Mux60~15 (
// Equation(s):
// \Mux60~15_combout  = (\Mux60~14_combout ) # ((!temp_imemload_output_16 & (\storeregister[2][3]~q  & temp_imemload_output_17)))

	.dataa(temp_imemload_output_16),
	.datab(\Mux60~14_combout ),
	.datac(\storeregister[2][3]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux60~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~15 .lut_mask = 16'hDCCC;
defparam \Mux60~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N22
cycloneive_lcell_comb \Mux60~16 (
// Equation(s):
// \Mux60~16_combout  = (temp_imemload_output_18 & ((\Mux60~13_combout ) # ((temp_imemload_output_19)))) # (!temp_imemload_output_18 & (((\Mux60~15_combout  & !temp_imemload_output_19))))

	.dataa(temp_imemload_output_18),
	.datab(\Mux60~13_combout ),
	.datac(\Mux60~15_combout ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux60~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~16 .lut_mask = 16'hAAD8;
defparam \Mux60~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N14
cycloneive_lcell_comb \Mux60~17 (
// Equation(s):
// \Mux60~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][3]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][3]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[12][3]~q ),
	.datad(\storeregister[13][3]~q ),
	.cin(gnd),
	.combout(\Mux60~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~17 .lut_mask = 16'hDC98;
defparam \Mux60~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N24
cycloneive_lcell_comb \Mux60~18 (
// Equation(s):
// \Mux60~18_combout  = (\Mux60~17_combout  & ((\storeregister[15][3]~q ) # ((!temp_imemload_output_17)))) # (!\Mux60~17_combout  & (((\storeregister[14][3]~q  & temp_imemload_output_17))))

	.dataa(\storeregister[15][3]~q ),
	.datab(\Mux60~17_combout ),
	.datac(\storeregister[14][3]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux60~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~18 .lut_mask = 16'hB8CC;
defparam \Mux60~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N4
cycloneive_lcell_comb \Mux60~10 (
// Equation(s):
// \Mux60~10_combout  = (temp_imemload_output_17 & ((temp_imemload_output_16) # ((\storeregister[10][3]~q )))) # (!temp_imemload_output_17 & (!temp_imemload_output_16 & ((\storeregister[8][3]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[10][3]~q ),
	.datad(\storeregister[8][3]~q ),
	.cin(gnd),
	.combout(\Mux60~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~10 .lut_mask = 16'hB9A8;
defparam \Mux60~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N8
cycloneive_lcell_comb \Mux60~11 (
// Equation(s):
// \Mux60~11_combout  = (\Mux60~10_combout  & ((\storeregister[11][3]~q ) # ((!temp_imemload_output_16)))) # (!\Mux60~10_combout  & (((\storeregister[9][3]~q  & temp_imemload_output_16))))

	.dataa(\storeregister[11][3]~q ),
	.datab(\storeregister[9][3]~q ),
	.datac(\Mux60~10_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux60~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~11 .lut_mask = 16'hACF0;
defparam \Mux60~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N8
cycloneive_lcell_comb \storeregister[29][16]~feeder (
// Equation(s):
// \storeregister[29][16]~feeder_combout  = Mux15

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux15),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[29][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][16]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[29][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N9
dffeas \storeregister[29][16] (
	.clk(!CLK),
	.d(\storeregister[29][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][16] .is_wysiwyg = "true";
defparam \storeregister[29][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N18
cycloneive_lcell_comb \storeregister[25][16]~feeder (
// Equation(s):
// \storeregister[25][16]~feeder_combout  = Mux15

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux15),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[25][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[25][16]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[25][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N19
dffeas \storeregister[25][16] (
	.clk(!CLK),
	.d(\storeregister[25][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][16] .is_wysiwyg = "true";
defparam \storeregister[25][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N17
dffeas \storeregister[17][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][16] .is_wysiwyg = "true";
defparam \storeregister[17][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N23
dffeas \storeregister[21][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][16] .is_wysiwyg = "true";
defparam \storeregister[21][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N22
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[21][16]~q ))) # (!temp_imemload_output_23 & (\storeregister[17][16]~q ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[17][16]~q ),
	.datac(\storeregister[21][16]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hFA44;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N30
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (temp_imemload_output_24 & ((\Mux15~0_combout  & (\storeregister[29][16]~q )) # (!\Mux15~0_combout  & ((\storeregister[25][16]~q ))))) # (!temp_imemload_output_24 & (((\Mux15~0_combout ))))

	.dataa(\storeregister[29][16]~q ),
	.datab(\storeregister[25][16]~q ),
	.datac(temp_imemload_output_24),
	.datad(\Mux15~0_combout ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hAFC0;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N6
cycloneive_lcell_comb \storeregister[26][16]~feeder (
// Equation(s):
// \storeregister[26][16]~feeder_combout  = Mux15

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux15),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[26][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[26][16]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[26][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N7
dffeas \storeregister[26][16] (
	.clk(!CLK),
	.d(\storeregister[26][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][16] .is_wysiwyg = "true";
defparam \storeregister[26][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N13
dffeas \storeregister[18][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][16] .is_wysiwyg = "true";
defparam \storeregister[18][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N12
cycloneive_lcell_comb \Mux15~2 (
// Equation(s):
// \Mux15~2_combout  = (temp_imemload_output_24 & ((\storeregister[26][16]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[18][16]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[26][16]~q ),
	.datac(\storeregister[18][16]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~2 .lut_mask = 16'hAAD8;
defparam \Mux15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N13
dffeas \storeregister[30][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][16] .is_wysiwyg = "true";
defparam \storeregister[30][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N10
cycloneive_lcell_comb \storeregister[22][16]~feeder (
// Equation(s):
// \storeregister[22][16]~feeder_combout  = Mux15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux15),
	.cin(gnd),
	.combout(\storeregister[22][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[22][16]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[22][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N11
dffeas \storeregister[22][16] (
	.clk(!CLK),
	.d(\storeregister[22][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][16] .is_wysiwyg = "true";
defparam \storeregister[22][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N16
cycloneive_lcell_comb \Mux15~3 (
// Equation(s):
// \Mux15~3_combout  = (temp_imemload_output_23 & ((\Mux15~2_combout  & (\storeregister[30][16]~q )) # (!\Mux15~2_combout  & ((\storeregister[22][16]~q ))))) # (!temp_imemload_output_23 & (\Mux15~2_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux15~2_combout ),
	.datac(\storeregister[30][16]~q ),
	.datad(\storeregister[22][16]~q ),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~3 .lut_mask = 16'hE6C4;
defparam \Mux15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N13
dffeas \storeregister[20][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][16] .is_wysiwyg = "true";
defparam \storeregister[20][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y35_N23
dffeas \storeregister[16][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][16] .is_wysiwyg = "true";
defparam \storeregister[16][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N30
cycloneive_lcell_comb \storeregister[24][16]~feeder (
// Equation(s):
// \storeregister[24][16]~feeder_combout  = Mux15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux15),
	.cin(gnd),
	.combout(\storeregister[24][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][16]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[24][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N31
dffeas \storeregister[24][16] (
	.clk(!CLK),
	.d(\storeregister[24][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][16] .is_wysiwyg = "true";
defparam \storeregister[24][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N22
cycloneive_lcell_comb \Mux15~4 (
// Equation(s):
// \Mux15~4_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[24][16]~q ))) # (!temp_imemload_output_24 & (\storeregister[16][16]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][16]~q ),
	.datad(\storeregister[24][16]~q ),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~4 .lut_mask = 16'hDC98;
defparam \Mux15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N2
cycloneive_lcell_comb \Mux15~5 (
// Equation(s):
// \Mux15~5_combout  = (temp_imemload_output_23 & ((\Mux15~4_combout  & (\storeregister[28][16]~q )) # (!\Mux15~4_combout  & ((\storeregister[20][16]~q ))))) # (!temp_imemload_output_23 & (((\Mux15~4_combout ))))

	.dataa(\storeregister[28][16]~q ),
	.datab(\storeregister[20][16]~q ),
	.datac(temp_imemload_output_23),
	.datad(\Mux15~4_combout ),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~5 .lut_mask = 16'hAFC0;
defparam \Mux15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N4
cycloneive_lcell_comb \Mux15~6 (
// Equation(s):
// \Mux15~6_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22)))) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\Mux15~3_combout )) # (!temp_imemload_output_22 & ((\Mux15~5_combout )))))

	.dataa(\Mux15~3_combout ),
	.datab(temp_imemload_output_21),
	.datac(temp_imemload_output_22),
	.datad(\Mux15~5_combout ),
	.cin(gnd),
	.combout(\Mux15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~6 .lut_mask = 16'hE3E0;
defparam \Mux15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N0
cycloneive_lcell_comb \storeregister[27][16]~feeder (
// Equation(s):
// \storeregister[27][16]~feeder_combout  = Mux15

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux15),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][16]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N1
dffeas \storeregister[27][16] (
	.clk(!CLK),
	.d(\storeregister[27][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][16] .is_wysiwyg = "true";
defparam \storeregister[27][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N13
dffeas \storeregister[23][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][16] .is_wysiwyg = "true";
defparam \storeregister[23][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N12
cycloneive_lcell_comb \Mux15~7 (
// Equation(s):
// \Mux15~7_combout  = (temp_imemload_output_23 & (((\storeregister[23][16]~q ) # (temp_imemload_output_24)))) # (!temp_imemload_output_23 & (\storeregister[19][16]~q  & ((!temp_imemload_output_24))))

	.dataa(\storeregister[19][16]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[23][16]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~7 .lut_mask = 16'hCCE2;
defparam \Mux15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N19
dffeas \storeregister[31][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][16] .is_wysiwyg = "true";
defparam \storeregister[31][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N16
cycloneive_lcell_comb \Mux15~8 (
// Equation(s):
// \Mux15~8_combout  = (temp_imemload_output_24 & ((\Mux15~7_combout  & ((\storeregister[31][16]~q ))) # (!\Mux15~7_combout  & (\storeregister[27][16]~q )))) # (!temp_imemload_output_24 & (((\Mux15~7_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[27][16]~q ),
	.datac(\Mux15~7_combout ),
	.datad(\storeregister[31][16]~q ),
	.cin(gnd),
	.combout(\Mux15~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~8 .lut_mask = 16'hF858;
defparam \Mux15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N1
dffeas \storeregister[10][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][16] .is_wysiwyg = "true";
defparam \storeregister[10][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N2
cycloneive_lcell_comb \storeregister[8][16]~feeder (
// Equation(s):
// \storeregister[8][16]~feeder_combout  = Mux15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux15),
	.cin(gnd),
	.combout(\storeregister[8][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[8][16]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[8][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N3
dffeas \storeregister[8][16] (
	.clk(!CLK),
	.d(\storeregister[8][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][16] .is_wysiwyg = "true";
defparam \storeregister[8][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N0
cycloneive_lcell_comb \Mux15~10 (
// Equation(s):
// \Mux15~10_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[10][16]~q )) # (!temp_imemload_output_22 & ((\storeregister[8][16]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][16]~q ),
	.datad(\storeregister[8][16]~q ),
	.cin(gnd),
	.combout(\Mux15~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~10 .lut_mask = 16'hD9C8;
defparam \Mux15~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N11
dffeas \storeregister[9][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][16] .is_wysiwyg = "true";
defparam \storeregister[9][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N29
dffeas \storeregister[11][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][16] .is_wysiwyg = "true";
defparam \storeregister[11][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N10
cycloneive_lcell_comb \Mux15~11 (
// Equation(s):
// \Mux15~11_combout  = (temp_imemload_output_21 & ((\Mux15~10_combout  & ((\storeregister[11][16]~q ))) # (!\Mux15~10_combout  & (\storeregister[9][16]~q )))) # (!temp_imemload_output_21 & (\Mux15~10_combout ))

	.dataa(temp_imemload_output_21),
	.datab(\Mux15~10_combout ),
	.datac(\storeregister[9][16]~q ),
	.datad(\storeregister[11][16]~q ),
	.cin(gnd),
	.combout(\Mux15~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~11 .lut_mask = 16'hEC64;
defparam \Mux15~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y40_N27
dffeas \storeregister[4][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][16] .is_wysiwyg = "true";
defparam \storeregister[4][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N25
dffeas \storeregister[5][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][16] .is_wysiwyg = "true";
defparam \storeregister[5][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N26
cycloneive_lcell_comb \Mux15~12 (
// Equation(s):
// \Mux15~12_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[5][16]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[4][16]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[4][16]~q ),
	.datad(\storeregister[5][16]~q ),
	.cin(gnd),
	.combout(\Mux15~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~12 .lut_mask = 16'hBA98;
defparam \Mux15~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N1
dffeas \storeregister[7][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][16] .is_wysiwyg = "true";
defparam \storeregister[7][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N0
cycloneive_lcell_comb \Mux15~13 (
// Equation(s):
// \Mux15~13_combout  = (\Mux15~12_combout  & (((\storeregister[7][16]~q ) # (!temp_imemload_output_22)))) # (!\Mux15~12_combout  & (\storeregister[6][16]~q  & ((temp_imemload_output_22))))

	.dataa(\storeregister[6][16]~q ),
	.datab(\Mux15~12_combout ),
	.datac(\storeregister[7][16]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux15~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~13 .lut_mask = 16'hE2CC;
defparam \Mux15~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N1
dffeas \storeregister[3][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][16] .is_wysiwyg = "true";
defparam \storeregister[3][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N7
dffeas \storeregister[1][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][16] .is_wysiwyg = "true";
defparam \storeregister[1][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N6
cycloneive_lcell_comb \Mux15~14 (
// Equation(s):
// \Mux15~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[3][16]~q )) # (!temp_imemload_output_22 & ((\storeregister[1][16]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[3][16]~q ),
	.datac(\storeregister[1][16]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux15~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~14 .lut_mask = 16'h88A0;
defparam \Mux15~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N30
cycloneive_lcell_comb \Mux15~15 (
// Equation(s):
// \Mux15~15_combout  = (\Mux15~14_combout ) # ((\storeregister[2][16]~q  & (!temp_imemload_output_21 & temp_imemload_output_22)))

	.dataa(\storeregister[2][16]~q ),
	.datab(temp_imemload_output_21),
	.datac(temp_imemload_output_22),
	.datad(\Mux15~14_combout ),
	.cin(gnd),
	.combout(\Mux15~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~15 .lut_mask = 16'hFF20;
defparam \Mux15~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N12
cycloneive_lcell_comb \Mux15~16 (
// Equation(s):
// \Mux15~16_combout  = (temp_imemload_output_23 & ((\Mux15~13_combout ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\Mux15~15_combout  & !temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\Mux15~13_combout ),
	.datac(\Mux15~15_combout ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux15~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~16 .lut_mask = 16'hAAD8;
defparam \Mux15~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N2
cycloneive_lcell_comb \storeregister[14][16]~feeder (
// Equation(s):
// \storeregister[14][16]~feeder_combout  = Mux15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux15),
	.cin(gnd),
	.combout(\storeregister[14][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][16]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N3
dffeas \storeregister[14][16] (
	.clk(!CLK),
	.d(\storeregister[14][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][16] .is_wysiwyg = "true";
defparam \storeregister[14][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N19
dffeas \storeregister[12][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][16] .is_wysiwyg = "true";
defparam \storeregister[12][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N9
dffeas \storeregister[13][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][16] .is_wysiwyg = "true";
defparam \storeregister[13][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N8
cycloneive_lcell_comb \Mux15~17 (
// Equation(s):
// \Mux15~17_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[13][16]~q ))) # (!temp_imemload_output_21 & (\storeregister[12][16]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[12][16]~q ),
	.datac(\storeregister[13][16]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux15~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~17 .lut_mask = 16'hFA44;
defparam \Mux15~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N20
cycloneive_lcell_comb \storeregister[15][16]~feeder (
// Equation(s):
// \storeregister[15][16]~feeder_combout  = Mux15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux15),
	.cin(gnd),
	.combout(\storeregister[15][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][16]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N21
dffeas \storeregister[15][16] (
	.clk(!CLK),
	.d(\storeregister[15][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][16] .is_wysiwyg = "true";
defparam \storeregister[15][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N6
cycloneive_lcell_comb \Mux15~18 (
// Equation(s):
// \Mux15~18_combout  = (temp_imemload_output_22 & ((\Mux15~17_combout  & ((\storeregister[15][16]~q ))) # (!\Mux15~17_combout  & (\storeregister[14][16]~q )))) # (!temp_imemload_output_22 & (((\Mux15~17_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[14][16]~q ),
	.datac(\Mux15~17_combout ),
	.datad(\storeregister[15][16]~q ),
	.cin(gnd),
	.combout(\Mux15~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~18 .lut_mask = 16'hF858;
defparam \Mux15~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N26
cycloneive_lcell_comb \storeregister[31][14]~feeder (
// Equation(s):
// \storeregister[31][14]~feeder_combout  = Mux17

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux17),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[31][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][14]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[31][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N27
dffeas \storeregister[31][14] (
	.clk(!CLK),
	.d(\storeregister[31][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][14] .is_wysiwyg = "true";
defparam \storeregister[31][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N29
dffeas \storeregister[27][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][14] .is_wysiwyg = "true";
defparam \storeregister[27][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N27
dffeas \storeregister[19][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][14] .is_wysiwyg = "true";
defparam \storeregister[19][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N5
dffeas \storeregister[23][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][14] .is_wysiwyg = "true";
defparam \storeregister[23][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N4
cycloneive_lcell_comb \Mux17~7 (
// Equation(s):
// \Mux17~7_combout  = (temp_imemload_output_23 & (((\storeregister[23][14]~q ) # (temp_imemload_output_24)))) # (!temp_imemload_output_23 & (\storeregister[19][14]~q  & ((!temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[19][14]~q ),
	.datac(\storeregister[23][14]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux17~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~7 .lut_mask = 16'hAAE4;
defparam \Mux17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N28
cycloneive_lcell_comb \Mux17~8 (
// Equation(s):
// \Mux17~8_combout  = (temp_imemload_output_24 & ((\Mux17~7_combout  & (\storeregister[31][14]~q )) # (!\Mux17~7_combout  & ((\storeregister[27][14]~q ))))) # (!temp_imemload_output_24 & (((\Mux17~7_combout ))))

	.dataa(\storeregister[31][14]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[27][14]~q ),
	.datad(\Mux17~7_combout ),
	.cin(gnd),
	.combout(\Mux17~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~8 .lut_mask = 16'hBBC0;
defparam \Mux17~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N5
dffeas \storeregister[30][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][14] .is_wysiwyg = "true";
defparam \storeregister[30][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N14
cycloneive_lcell_comb \storeregister[26][14]~feeder (
// Equation(s):
// \storeregister[26][14]~feeder_combout  = Mux17

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux17),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[26][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[26][14]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[26][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N15
dffeas \storeregister[26][14] (
	.clk(!CLK),
	.d(\storeregister[26][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][14] .is_wysiwyg = "true";
defparam \storeregister[26][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N29
dffeas \storeregister[18][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][14] .is_wysiwyg = "true";
defparam \storeregister[18][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N28
cycloneive_lcell_comb \Mux17~2 (
// Equation(s):
// \Mux17~2_combout  = (temp_imemload_output_24 & ((\storeregister[26][14]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[18][14]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[26][14]~q ),
	.datac(\storeregister[18][14]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~2 .lut_mask = 16'hAAD8;
defparam \Mux17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N19
dffeas \storeregister[22][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][14] .is_wysiwyg = "true";
defparam \storeregister[22][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N28
cycloneive_lcell_comb \Mux17~3 (
// Equation(s):
// \Mux17~3_combout  = (temp_imemload_output_23 & ((\Mux17~2_combout  & (\storeregister[30][14]~q )) # (!\Mux17~2_combout  & ((\storeregister[22][14]~q ))))) # (!temp_imemload_output_23 & (((\Mux17~2_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[30][14]~q ),
	.datac(\Mux17~2_combout ),
	.datad(\storeregister[22][14]~q ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~3 .lut_mask = 16'hDAD0;
defparam \Mux17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N17
dffeas \storeregister[16][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][14] .is_wysiwyg = "true";
defparam \storeregister[16][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N11
dffeas \storeregister[24][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][14] .is_wysiwyg = "true";
defparam \storeregister[24][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N10
cycloneive_lcell_comb \Mux17~4 (
// Equation(s):
// \Mux17~4_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[24][14]~q ))) # (!temp_imemload_output_24 & (\storeregister[16][14]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[16][14]~q ),
	.datac(\storeregister[24][14]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~4 .lut_mask = 16'hFA44;
defparam \Mux17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N7
dffeas \storeregister[20][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][14] .is_wysiwyg = "true";
defparam \storeregister[20][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N13
dffeas \storeregister[28][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][14] .is_wysiwyg = "true";
defparam \storeregister[28][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N6
cycloneive_lcell_comb \Mux17~5 (
// Equation(s):
// \Mux17~5_combout  = (temp_imemload_output_23 & ((\Mux17~4_combout  & ((\storeregister[28][14]~q ))) # (!\Mux17~4_combout  & (\storeregister[20][14]~q )))) # (!temp_imemload_output_23 & (\Mux17~4_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux17~4_combout ),
	.datac(\storeregister[20][14]~q ),
	.datad(\storeregister[28][14]~q ),
	.cin(gnd),
	.combout(\Mux17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~5 .lut_mask = 16'hEC64;
defparam \Mux17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N24
cycloneive_lcell_comb \Mux17~6 (
// Equation(s):
// \Mux17~6_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\Mux17~3_combout )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & ((\Mux17~5_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\Mux17~3_combout ),
	.datad(\Mux17~5_combout ),
	.cin(gnd),
	.combout(\Mux17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~6 .lut_mask = 16'hB9A8;
defparam \Mux17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N22
cycloneive_lcell_comb \storeregister[29][14]~feeder (
// Equation(s):
// \storeregister[29][14]~feeder_combout  = Mux17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux17),
	.cin(gnd),
	.combout(\storeregister[29][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][14]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[29][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N23
dffeas \storeregister[29][14] (
	.clk(!CLK),
	.d(\storeregister[29][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][14] .is_wysiwyg = "true";
defparam \storeregister[29][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N30
cycloneive_lcell_comb \storeregister[25][14]~feeder (
// Equation(s):
// \storeregister[25][14]~feeder_combout  = Mux17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux17),
	.cin(gnd),
	.combout(\storeregister[25][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[25][14]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[25][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N31
dffeas \storeregister[25][14] (
	.clk(!CLK),
	.d(\storeregister[25][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][14] .is_wysiwyg = "true";
defparam \storeregister[25][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N28
cycloneive_lcell_comb \storeregister[21][14]~feeder (
// Equation(s):
// \storeregister[21][14]~feeder_combout  = Mux17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux17),
	.cin(gnd),
	.combout(\storeregister[21][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][14]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[21][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N29
dffeas \storeregister[21][14] (
	.clk(!CLK),
	.d(\storeregister[21][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][14] .is_wysiwyg = "true";
defparam \storeregister[21][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N23
dffeas \storeregister[17][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][14] .is_wysiwyg = "true";
defparam \storeregister[17][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N22
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (temp_imemload_output_23 & ((\storeregister[21][14]~q ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\storeregister[17][14]~q  & !temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[21][14]~q ),
	.datac(\storeregister[17][14]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hAAD8;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N20
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (temp_imemload_output_24 & ((\Mux17~0_combout  & (\storeregister[29][14]~q )) # (!\Mux17~0_combout  & ((\storeregister[25][14]~q ))))) # (!temp_imemload_output_24 & (((\Mux17~0_combout ))))

	.dataa(\storeregister[29][14]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[25][14]~q ),
	.datad(\Mux17~0_combout ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hBBC0;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N19
dffeas \storeregister[12][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][14] .is_wysiwyg = "true";
defparam \storeregister[12][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N26
cycloneive_lcell_comb \storeregister[13][14]~feeder (
// Equation(s):
// \storeregister[13][14]~feeder_combout  = Mux17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux17),
	.cin(gnd),
	.combout(\storeregister[13][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[13][14]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[13][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N27
dffeas \storeregister[13][14] (
	.clk(!CLK),
	.d(\storeregister[13][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][14] .is_wysiwyg = "true";
defparam \storeregister[13][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N20
cycloneive_lcell_comb \Mux17~17 (
// Equation(s):
// \Mux17~17_combout  = (temp_imemload_output_21 & (((\storeregister[13][14]~q ) # (temp_imemload_output_22)))) # (!temp_imemload_output_21 & (\storeregister[12][14]~q  & ((!temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[12][14]~q ),
	.datac(\storeregister[13][14]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux17~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~17 .lut_mask = 16'hAAE4;
defparam \Mux17~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N4
cycloneive_lcell_comb \storeregister[15][14]~feeder (
// Equation(s):
// \storeregister[15][14]~feeder_combout  = Mux17

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux17),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[15][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][14]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[15][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N5
dffeas \storeregister[15][14] (
	.clk(!CLK),
	.d(\storeregister[15][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][14] .is_wysiwyg = "true";
defparam \storeregister[15][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N2
cycloneive_lcell_comb \storeregister[14][14]~feeder (
// Equation(s):
// \storeregister[14][14]~feeder_combout  = Mux17

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux17),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[14][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][14]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[14][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N3
dffeas \storeregister[14][14] (
	.clk(!CLK),
	.d(\storeregister[14][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][14] .is_wysiwyg = "true";
defparam \storeregister[14][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N6
cycloneive_lcell_comb \Mux17~18 (
// Equation(s):
// \Mux17~18_combout  = (\Mux17~17_combout  & (((\storeregister[15][14]~q )) # (!temp_imemload_output_22))) # (!\Mux17~17_combout  & (temp_imemload_output_22 & ((\storeregister[14][14]~q ))))

	.dataa(\Mux17~17_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[15][14]~q ),
	.datad(\storeregister[14][14]~q ),
	.cin(gnd),
	.combout(\Mux17~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~18 .lut_mask = 16'hE6A2;
defparam \Mux17~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N9
dffeas \storeregister[9][14] (
	.clk(!CLK),
	.d(Mux17),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][14] .is_wysiwyg = "true";
defparam \storeregister[9][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N31
dffeas \storeregister[10][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][14] .is_wysiwyg = "true";
defparam \storeregister[10][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N8
cycloneive_lcell_comb \storeregister[8][14]~feeder (
// Equation(s):
// \storeregister[8][14]~feeder_combout  = Mux17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux17),
	.cin(gnd),
	.combout(\storeregister[8][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[8][14]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[8][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N9
dffeas \storeregister[8][14] (
	.clk(!CLK),
	.d(\storeregister[8][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][14] .is_wysiwyg = "true";
defparam \storeregister[8][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N30
cycloneive_lcell_comb \Mux17~10 (
// Equation(s):
// \Mux17~10_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[10][14]~q )) # (!temp_imemload_output_22 & ((\storeregister[8][14]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][14]~q ),
	.datad(\storeregister[8][14]~q ),
	.cin(gnd),
	.combout(\Mux17~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~10 .lut_mask = 16'hD9C8;
defparam \Mux17~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N17
dffeas \storeregister[11][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][14] .is_wysiwyg = "true";
defparam \storeregister[11][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N0
cycloneive_lcell_comb \Mux17~11 (
// Equation(s):
// \Mux17~11_combout  = (temp_imemload_output_21 & ((\Mux17~10_combout  & ((\storeregister[11][14]~q ))) # (!\Mux17~10_combout  & (\storeregister[9][14]~q )))) # (!temp_imemload_output_21 & (((\Mux17~10_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[9][14]~q ),
	.datac(\Mux17~10_combout ),
	.datad(\storeregister[11][14]~q ),
	.cin(gnd),
	.combout(\Mux17~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~11 .lut_mask = 16'hF858;
defparam \Mux17~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N19
dffeas \storeregister[6][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][14] .is_wysiwyg = "true";
defparam \storeregister[6][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N13
dffeas \storeregister[7][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][14] .is_wysiwyg = "true";
defparam \storeregister[7][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N12
cycloneive_lcell_comb \Mux17~13 (
// Equation(s):
// \Mux17~13_combout  = (\Mux17~12_combout  & (((\storeregister[7][14]~q ) # (!temp_imemload_output_22)))) # (!\Mux17~12_combout  & (\storeregister[6][14]~q  & ((temp_imemload_output_22))))

	.dataa(\Mux17~12_combout ),
	.datab(\storeregister[6][14]~q ),
	.datac(\storeregister[7][14]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux17~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~13 .lut_mask = 16'hE4AA;
defparam \Mux17~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N15
dffeas \storeregister[2][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][14] .is_wysiwyg = "true";
defparam \storeregister[2][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N18
cycloneive_lcell_comb \Mux17~15 (
// Equation(s):
// \Mux17~15_combout  = (\Mux17~14_combout ) # ((temp_imemload_output_22 & (\storeregister[2][14]~q  & !temp_imemload_output_21)))

	.dataa(\Mux17~14_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][14]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux17~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~15 .lut_mask = 16'hAAEA;
defparam \Mux17~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N0
cycloneive_lcell_comb \Mux17~16 (
// Equation(s):
// \Mux17~16_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\Mux17~13_combout )) # (!temp_imemload_output_23 & ((\Mux17~15_combout )))))

	.dataa(\Mux17~13_combout ),
	.datab(temp_imemload_output_24),
	.datac(temp_imemload_output_23),
	.datad(\Mux17~15_combout ),
	.cin(gnd),
	.combout(\Mux17~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~16 .lut_mask = 16'hE3E0;
defparam \Mux17~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N1
dffeas \storeregister[28][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][15] .is_wysiwyg = "true";
defparam \storeregister[28][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N27
dffeas \storeregister[24][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][15] .is_wysiwyg = "true";
defparam \storeregister[24][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N26
cycloneive_lcell_comb \Mux16~5 (
// Equation(s):
// \Mux16~5_combout  = (\Mux16~4_combout  & ((\storeregister[28][15]~q ) # ((!temp_imemload_output_24)))) # (!\Mux16~4_combout  & (((\storeregister[24][15]~q  & temp_imemload_output_24))))

	.dataa(\Mux16~4_combout ),
	.datab(\storeregister[28][15]~q ),
	.datac(\storeregister[24][15]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~5 .lut_mask = 16'hD8AA;
defparam \Mux16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N9
dffeas \storeregister[22][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][15] .is_wysiwyg = "true";
defparam \storeregister[22][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N15
dffeas \storeregister[18][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][15] .is_wysiwyg = "true";
defparam \storeregister[18][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N8
cycloneive_lcell_comb \Mux16~2 (
// Equation(s):
// \Mux16~2_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[22][15]~q )) # (!temp_imemload_output_23 & ((\storeregister[18][15]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[22][15]~q ),
	.datad(\storeregister[18][15]~q ),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~2 .lut_mask = 16'hD9C8;
defparam \Mux16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N27
dffeas \storeregister[30][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][15] .is_wysiwyg = "true";
defparam \storeregister[30][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N30
cycloneive_lcell_comb \storeregister[26][15]~feeder (
// Equation(s):
// \storeregister[26][15]~feeder_combout  = Mux16

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux16),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[26][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[26][15]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[26][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N31
dffeas \storeregister[26][15] (
	.clk(!CLK),
	.d(\storeregister[26][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][15] .is_wysiwyg = "true";
defparam \storeregister[26][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N26
cycloneive_lcell_comb \Mux16~3 (
// Equation(s):
// \Mux16~3_combout  = (temp_imemload_output_24 & ((\Mux16~2_combout  & (\storeregister[30][15]~q )) # (!\Mux16~2_combout  & ((\storeregister[26][15]~q ))))) # (!temp_imemload_output_24 & (\Mux16~2_combout ))

	.dataa(temp_imemload_output_24),
	.datab(\Mux16~2_combout ),
	.datac(\storeregister[30][15]~q ),
	.datad(\storeregister[26][15]~q ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~3 .lut_mask = 16'hE6C4;
defparam \Mux16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N22
cycloneive_lcell_comb \Mux16~6 (
// Equation(s):
// \Mux16~6_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\Mux16~3_combout )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & (\Mux16~5_combout )))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\Mux16~5_combout ),
	.datad(\Mux16~3_combout ),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~6 .lut_mask = 16'hBA98;
defparam \Mux16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N20
cycloneive_lcell_comb \storeregister[29][15]~feeder (
// Equation(s):
// \storeregister[29][15]~feeder_combout  = Mux16

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux16),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[29][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][15]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[29][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N21
dffeas \storeregister[29][15] (
	.clk(!CLK),
	.d(\storeregister[29][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][15] .is_wysiwyg = "true";
defparam \storeregister[29][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N25
dffeas \storeregister[21][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][15] .is_wysiwyg = "true";
defparam \storeregister[21][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N24
cycloneive_lcell_comb \storeregister[25][15]~feeder (
// Equation(s):
// \storeregister[25][15]~feeder_combout  = Mux16

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux16),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[25][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[25][15]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[25][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N25
dffeas \storeregister[25][15] (
	.clk(!CLK),
	.d(\storeregister[25][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][15] .is_wysiwyg = "true";
defparam \storeregister[25][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N19
dffeas \storeregister[17][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][15] .is_wysiwyg = "true";
defparam \storeregister[17][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N18
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (temp_imemload_output_24 & ((\storeregister[25][15]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[17][15]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[25][15]~q ),
	.datac(\storeregister[17][15]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hAAD8;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N4
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (temp_imemload_output_23 & ((\Mux16~0_combout  & (\storeregister[29][15]~q )) # (!\Mux16~0_combout  & ((\storeregister[21][15]~q ))))) # (!temp_imemload_output_23 & (((\Mux16~0_combout ))))

	.dataa(\storeregister[29][15]~q ),
	.datab(\storeregister[21][15]~q ),
	.datac(temp_imemload_output_23),
	.datad(\Mux16~0_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hAFC0;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N1
dffeas \storeregister[27][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][15] .is_wysiwyg = "true";
defparam \storeregister[27][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N0
cycloneive_lcell_comb \Mux16~7 (
// Equation(s):
// \Mux16~7_combout  = (temp_imemload_output_24 & (((\storeregister[27][15]~q ) # (temp_imemload_output_23)))) # (!temp_imemload_output_24 & (\storeregister[19][15]~q  & ((!temp_imemload_output_23))))

	.dataa(\storeregister[19][15]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[27][15]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~7 .lut_mask = 16'hCCE2;
defparam \Mux16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N14
cycloneive_lcell_comb \storeregister[23][15]~feeder (
// Equation(s):
// \storeregister[23][15]~feeder_combout  = Mux16

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux16),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[23][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][15]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[23][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N15
dffeas \storeregister[23][15] (
	.clk(!CLK),
	.d(\storeregister[23][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][15] .is_wysiwyg = "true";
defparam \storeregister[23][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N28
cycloneive_lcell_comb \storeregister[31][15]~feeder (
// Equation(s):
// \storeregister[31][15]~feeder_combout  = Mux16

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux16),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[31][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][15]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[31][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N29
dffeas \storeregister[31][15] (
	.clk(!CLK),
	.d(\storeregister[31][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][15] .is_wysiwyg = "true";
defparam \storeregister[31][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N4
cycloneive_lcell_comb \Mux16~8 (
// Equation(s):
// \Mux16~8_combout  = (temp_imemload_output_23 & ((\Mux16~7_combout  & ((\storeregister[31][15]~q ))) # (!\Mux16~7_combout  & (\storeregister[23][15]~q )))) # (!temp_imemload_output_23 & (\Mux16~7_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux16~7_combout ),
	.datac(\storeregister[23][15]~q ),
	.datad(\storeregister[31][15]~q ),
	.cin(gnd),
	.combout(\Mux16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~8 .lut_mask = 16'hEC64;
defparam \Mux16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N23
dffeas \storeregister[7][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][15] .is_wysiwyg = "true";
defparam \storeregister[7][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N25
dffeas \storeregister[6][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][15] .is_wysiwyg = "true";
defparam \storeregister[6][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y42_N3
dffeas \storeregister[4][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][15] .is_wysiwyg = "true";
defparam \storeregister[4][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y42_N25
dffeas \storeregister[5][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][15] .is_wysiwyg = "true";
defparam \storeregister[5][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N24
cycloneive_lcell_comb \Mux16~10 (
// Equation(s):
// \Mux16~10_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[5][15]~q ))) # (!temp_imemload_output_21 & (\storeregister[4][15]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[4][15]~q ),
	.datac(\storeregister[5][15]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~10 .lut_mask = 16'hFA44;
defparam \Mux16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N24
cycloneive_lcell_comb \Mux16~11 (
// Equation(s):
// \Mux16~11_combout  = (temp_imemload_output_22 & ((\Mux16~10_combout  & (\storeregister[7][15]~q )) # (!\Mux16~10_combout  & ((\storeregister[6][15]~q ))))) # (!temp_imemload_output_22 & (((\Mux16~10_combout ))))

	.dataa(\storeregister[7][15]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[6][15]~q ),
	.datad(\Mux16~10_combout ),
	.cin(gnd),
	.combout(\Mux16~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~11 .lut_mask = 16'hBBC0;
defparam \Mux16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N28
cycloneive_lcell_comb \storeregister[15][15]~feeder (
// Equation(s):
// \storeregister[15][15]~feeder_combout  = Mux16

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux16),
	.cin(gnd),
	.combout(\storeregister[15][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][15]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N29
dffeas \storeregister[15][15] (
	.clk(!CLK),
	.d(\storeregister[15][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][15] .is_wysiwyg = "true";
defparam \storeregister[15][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N27
dffeas \storeregister[12][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][15] .is_wysiwyg = "true";
defparam \storeregister[12][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N17
dffeas \storeregister[13][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][15] .is_wysiwyg = "true";
defparam \storeregister[13][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N16
cycloneive_lcell_comb \Mux16~17 (
// Equation(s):
// \Mux16~17_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[13][15]~q ))) # (!temp_imemload_output_21 & (\storeregister[12][15]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[12][15]~q ),
	.datac(\storeregister[13][15]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux16~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~17 .lut_mask = 16'hFA44;
defparam \Mux16~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N18
cycloneive_lcell_comb \storeregister[14][15]~feeder (
// Equation(s):
// \storeregister[14][15]~feeder_combout  = Mux16

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux16),
	.cin(gnd),
	.combout(\storeregister[14][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][15]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N19
dffeas \storeregister[14][15] (
	.clk(!CLK),
	.d(\storeregister[14][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][15] .is_wysiwyg = "true";
defparam \storeregister[14][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N22
cycloneive_lcell_comb \Mux16~18 (
// Equation(s):
// \Mux16~18_combout  = (temp_imemload_output_22 & ((\Mux16~17_combout  & (\storeregister[15][15]~q )) # (!\Mux16~17_combout  & ((\storeregister[14][15]~q ))))) # (!temp_imemload_output_22 & (((\Mux16~17_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[15][15]~q ),
	.datac(\Mux16~17_combout ),
	.datad(\storeregister[14][15]~q ),
	.cin(gnd),
	.combout(\Mux16~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~18 .lut_mask = 16'hDAD0;
defparam \Mux16~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N9
dffeas \storeregister[3][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][15] .is_wysiwyg = "true";
defparam \storeregister[3][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N11
dffeas \storeregister[1][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][15] .is_wysiwyg = "true";
defparam \storeregister[1][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N10
cycloneive_lcell_comb \Mux16~14 (
// Equation(s):
// \Mux16~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[3][15]~q )) # (!temp_imemload_output_22 & ((\storeregister[1][15]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[3][15]~q ),
	.datac(\storeregister[1][15]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux16~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~14 .lut_mask = 16'h88A0;
defparam \Mux16~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N21
dffeas \storeregister[2][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][15] .is_wysiwyg = "true";
defparam \storeregister[2][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N10
cycloneive_lcell_comb \Mux16~15 (
// Equation(s):
// \Mux16~15_combout  = (\Mux16~14_combout ) # ((temp_imemload_output_22 & (!temp_imemload_output_21 & \storeregister[2][15]~q )))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\Mux16~14_combout ),
	.datad(\storeregister[2][15]~q ),
	.cin(gnd),
	.combout(\Mux16~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~15 .lut_mask = 16'hF2F0;
defparam \Mux16~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N31
dffeas \storeregister[11][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][15] .is_wysiwyg = "true";
defparam \storeregister[11][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N1
dffeas \storeregister[9][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][15] .is_wysiwyg = "true";
defparam \storeregister[9][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N30
cycloneive_lcell_comb \Mux16~13 (
// Equation(s):
// \Mux16~13_combout  = (\Mux16~12_combout  & (((\storeregister[11][15]~q )) # (!temp_imemload_output_21))) # (!\Mux16~12_combout  & (temp_imemload_output_21 & ((\storeregister[9][15]~q ))))

	.dataa(\Mux16~12_combout ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[11][15]~q ),
	.datad(\storeregister[9][15]~q ),
	.cin(gnd),
	.combout(\Mux16~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~13 .lut_mask = 16'hE6A2;
defparam \Mux16~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N18
cycloneive_lcell_comb \Mux16~16 (
// Equation(s):
// \Mux16~16_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23) # (\Mux16~13_combout )))) # (!temp_imemload_output_24 & (\Mux16~15_combout  & (!temp_imemload_output_23)))

	.dataa(\Mux16~15_combout ),
	.datab(temp_imemload_output_24),
	.datac(temp_imemload_output_23),
	.datad(\Mux16~13_combout ),
	.cin(gnd),
	.combout(\Mux16~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~16 .lut_mask = 16'hCEC2;
defparam \Mux16~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N17
dffeas \storeregister[23][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][13] .is_wysiwyg = "true";
defparam \storeregister[23][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N21
dffeas \storeregister[27][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][13] .is_wysiwyg = "true";
defparam \storeregister[27][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N17
dffeas \storeregister[19][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][13] .is_wysiwyg = "true";
defparam \storeregister[19][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N16
cycloneive_lcell_comb \Mux18~7 (
// Equation(s):
// \Mux18~7_combout  = (temp_imemload_output_24 & ((\storeregister[27][13]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[19][13]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[27][13]~q ),
	.datac(\storeregister[19][13]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~7 .lut_mask = 16'hAAD8;
defparam \Mux18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N19
dffeas \storeregister[31][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][13] .is_wysiwyg = "true";
defparam \storeregister[31][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N18
cycloneive_lcell_comb \Mux18~8 (
// Equation(s):
// \Mux18~8_combout  = (\Mux18~7_combout  & (((\storeregister[31][13]~q ) # (!temp_imemload_output_23)))) # (!\Mux18~7_combout  & (\storeregister[23][13]~q  & ((temp_imemload_output_23))))

	.dataa(\storeregister[23][13]~q ),
	.datab(\Mux18~7_combout ),
	.datac(\storeregister[31][13]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux18~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~8 .lut_mask = 16'hE2CC;
defparam \Mux18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N17
dffeas \storeregister[25][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][13] .is_wysiwyg = "true";
defparam \storeregister[25][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N16
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (temp_imemload_output_24 & (((\storeregister[25][13]~q ) # (temp_imemload_output_23)))) # (!temp_imemload_output_24 & (\storeregister[17][13]~q  & ((!temp_imemload_output_23))))

	.dataa(\storeregister[17][13]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[25][13]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hCCE2;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N2
cycloneive_lcell_comb \storeregister[21][13]~feeder (
// Equation(s):
// \storeregister[21][13]~feeder_combout  = Mux18

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux18),
	.cin(gnd),
	.combout(\storeregister[21][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][13]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[21][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N3
dffeas \storeregister[21][13] (
	.clk(!CLK),
	.d(\storeregister[21][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][13] .is_wysiwyg = "true";
defparam \storeregister[21][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N2
cycloneive_lcell_comb \storeregister[29][13]~feeder (
// Equation(s):
// \storeregister[29][13]~feeder_combout  = Mux18

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux18),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[29][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][13]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[29][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N3
dffeas \storeregister[29][13] (
	.clk(!CLK),
	.d(\storeregister[29][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][13] .is_wysiwyg = "true";
defparam \storeregister[29][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N28
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (temp_imemload_output_23 & ((\Mux18~0_combout  & ((\storeregister[29][13]~q ))) # (!\Mux18~0_combout  & (\storeregister[21][13]~q )))) # (!temp_imemload_output_23 & (\Mux18~0_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux18~0_combout ),
	.datac(\storeregister[21][13]~q ),
	.datad(\storeregister[29][13]~q ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hEC64;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N17
dffeas \storeregister[22][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][13] .is_wysiwyg = "true";
defparam \storeregister[22][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N31
dffeas \storeregister[18][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][13] .is_wysiwyg = "true";
defparam \storeregister[18][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N30
cycloneive_lcell_comb \Mux18~2 (
// Equation(s):
// \Mux18~2_combout  = (temp_imemload_output_23 & ((\storeregister[22][13]~q ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\storeregister[18][13]~q  & !temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[22][13]~q ),
	.datac(\storeregister[18][13]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~2 .lut_mask = 16'hAAD8;
defparam \Mux18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N7
dffeas \storeregister[30][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][13] .is_wysiwyg = "true";
defparam \storeregister[30][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N13
dffeas \storeregister[26][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][13] .is_wysiwyg = "true";
defparam \storeregister[26][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N6
cycloneive_lcell_comb \Mux18~3 (
// Equation(s):
// \Mux18~3_combout  = (temp_imemload_output_24 & ((\Mux18~2_combout  & (\storeregister[30][13]~q )) # (!\Mux18~2_combout  & ((\storeregister[26][13]~q ))))) # (!temp_imemload_output_24 & (\Mux18~2_combout ))

	.dataa(temp_imemload_output_24),
	.datab(\Mux18~2_combout ),
	.datac(\storeregister[30][13]~q ),
	.datad(\storeregister[26][13]~q ),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~3 .lut_mask = 16'hE6C4;
defparam \Mux18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N19
dffeas \storeregister[24][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][13] .is_wysiwyg = "true";
defparam \storeregister[24][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N28
cycloneive_lcell_comb \storeregister[28][13]~feeder (
// Equation(s):
// \storeregister[28][13]~feeder_combout  = Mux18

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux18),
	.cin(gnd),
	.combout(\storeregister[28][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][13]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[28][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N29
dffeas \storeregister[28][13] (
	.clk(!CLK),
	.d(\storeregister[28][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][13] .is_wysiwyg = "true";
defparam \storeregister[28][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N22
cycloneive_lcell_comb \Mux18~5 (
// Equation(s):
// \Mux18~5_combout  = (\Mux18~4_combout  & (((\storeregister[28][13]~q ) # (!temp_imemload_output_24)))) # (!\Mux18~4_combout  & (\storeregister[24][13]~q  & (temp_imemload_output_24)))

	.dataa(\Mux18~4_combout ),
	.datab(\storeregister[24][13]~q ),
	.datac(temp_imemload_output_24),
	.datad(\storeregister[28][13]~q ),
	.cin(gnd),
	.combout(\Mux18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~5 .lut_mask = 16'hEA4A;
defparam \Mux18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N24
cycloneive_lcell_comb \Mux18~6 (
// Equation(s):
// \Mux18~6_combout  = (temp_imemload_output_22 & ((\Mux18~3_combout ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((\Mux18~5_combout  & !temp_imemload_output_21))))

	.dataa(temp_imemload_output_22),
	.datab(\Mux18~3_combout ),
	.datac(\Mux18~5_combout ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~6 .lut_mask = 16'hAAD8;
defparam \Mux18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N27
dffeas \storeregister[11][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][13] .is_wysiwyg = "true";
defparam \storeregister[11][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N13
dffeas \storeregister[9][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][13] .is_wysiwyg = "true";
defparam \storeregister[9][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N26
cycloneive_lcell_comb \Mux18~13 (
// Equation(s):
// \Mux18~13_combout  = (\Mux18~12_combout  & (((\storeregister[11][13]~q )) # (!temp_imemload_output_21))) # (!\Mux18~12_combout  & (temp_imemload_output_21 & ((\storeregister[9][13]~q ))))

	.dataa(\Mux18~12_combout ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[11][13]~q ),
	.datad(\storeregister[9][13]~q ),
	.cin(gnd),
	.combout(\Mux18~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~13 .lut_mask = 16'hE6A2;
defparam \Mux18~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N8
cycloneive_lcell_comb \storeregister[2][13]~feeder (
// Equation(s):
// \storeregister[2][13]~feeder_combout  = Mux18

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux18),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[2][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[2][13]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[2][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N9
dffeas \storeregister[2][13] (
	.clk(!CLK),
	.d(\storeregister[2][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][13] .is_wysiwyg = "true";
defparam \storeregister[2][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N23
dffeas \storeregister[1][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][13] .is_wysiwyg = "true";
defparam \storeregister[1][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N21
dffeas \storeregister[3][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][13] .is_wysiwyg = "true";
defparam \storeregister[3][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N20
cycloneive_lcell_comb \Mux18~14 (
// Equation(s):
// \Mux18~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][13]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][13]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[1][13]~q ),
	.datac(\storeregister[3][13]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux18~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~14 .lut_mask = 16'hA088;
defparam \Mux18~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N14
cycloneive_lcell_comb \Mux18~15 (
// Equation(s):
// \Mux18~15_combout  = (\Mux18~14_combout ) # ((!temp_imemload_output_21 & (\storeregister[2][13]~q  & temp_imemload_output_22)))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[2][13]~q ),
	.datac(temp_imemload_output_22),
	.datad(\Mux18~14_combout ),
	.cin(gnd),
	.combout(\Mux18~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~15 .lut_mask = 16'hFF40;
defparam \Mux18~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N30
cycloneive_lcell_comb \Mux18~16 (
// Equation(s):
// \Mux18~16_combout  = (temp_imemload_output_24 & ((\Mux18~13_combout ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((!temp_imemload_output_23 & \Mux18~15_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\Mux18~13_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux18~15_combout ),
	.cin(gnd),
	.combout(\Mux18~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~16 .lut_mask = 16'hADA8;
defparam \Mux18~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N7
dffeas \storeregister[7][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][13] .is_wysiwyg = "true";
defparam \storeregister[7][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N1
dffeas \storeregister[6][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][13] .is_wysiwyg = "true";
defparam \storeregister[6][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y41_N29
dffeas \storeregister[5][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][13] .is_wysiwyg = "true";
defparam \storeregister[5][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N28
cycloneive_lcell_comb \Mux18~10 (
// Equation(s):
// \Mux18~10_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[5][13]~q ))) # (!temp_imemload_output_21 & (\storeregister[4][13]~q ))))

	.dataa(\storeregister[4][13]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[5][13]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux18~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~10 .lut_mask = 16'hFC22;
defparam \Mux18~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N0
cycloneive_lcell_comb \Mux18~11 (
// Equation(s):
// \Mux18~11_combout  = (temp_imemload_output_22 & ((\Mux18~10_combout  & (\storeregister[7][13]~q )) # (!\Mux18~10_combout  & ((\storeregister[6][13]~q ))))) # (!temp_imemload_output_22 & (((\Mux18~10_combout ))))

	.dataa(\storeregister[7][13]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[6][13]~q ),
	.datad(\Mux18~10_combout ),
	.cin(gnd),
	.combout(\Mux18~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~11 .lut_mask = 16'hBBC0;
defparam \Mux18~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N26
cycloneive_lcell_comb \storeregister[14][13]~feeder (
// Equation(s):
// \storeregister[14][13]~feeder_combout  = Mux18

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux18),
	.cin(gnd),
	.combout(\storeregister[14][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][13]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N27
dffeas \storeregister[14][13] (
	.clk(!CLK),
	.d(\storeregister[14][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][13] .is_wysiwyg = "true";
defparam \storeregister[14][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N9
dffeas \storeregister[13][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][13] .is_wysiwyg = "true";
defparam \storeregister[13][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N23
dffeas \storeregister[12][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][13] .is_wysiwyg = "true";
defparam \storeregister[12][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N22
cycloneive_lcell_comb \Mux18~17 (
// Equation(s):
// \Mux18~17_combout  = (temp_imemload_output_21 & ((\storeregister[13][13]~q ) # ((temp_imemload_output_22)))) # (!temp_imemload_output_21 & (((\storeregister[12][13]~q  & !temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[13][13]~q ),
	.datac(\storeregister[12][13]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux18~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~17 .lut_mask = 16'hAAD8;
defparam \Mux18~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N0
cycloneive_lcell_comb \storeregister[15][13]~feeder (
// Equation(s):
// \storeregister[15][13]~feeder_combout  = Mux18

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux18),
	.cin(gnd),
	.combout(\storeregister[15][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][13]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N1
dffeas \storeregister[15][13] (
	.clk(!CLK),
	.d(\storeregister[15][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][13] .is_wysiwyg = "true";
defparam \storeregister[15][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N18
cycloneive_lcell_comb \Mux18~18 (
// Equation(s):
// \Mux18~18_combout  = (\Mux18~17_combout  & (((\storeregister[15][13]~q ) # (!temp_imemload_output_22)))) # (!\Mux18~17_combout  & (\storeregister[14][13]~q  & (temp_imemload_output_22)))

	.dataa(\storeregister[14][13]~q ),
	.datab(\Mux18~17_combout ),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[15][13]~q ),
	.cin(gnd),
	.combout(\Mux18~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~18 .lut_mask = 16'hEC2C;
defparam \Mux18~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N18
cycloneive_lcell_comb \storeregister[29][12]~feeder (
// Equation(s):
// \storeregister[29][12]~feeder_combout  = Mux19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux19),
	.cin(gnd),
	.combout(\storeregister[29][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][12]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[29][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N19
dffeas \storeregister[29][12] (
	.clk(!CLK),
	.d(\storeregister[29][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][12] .is_wysiwyg = "true";
defparam \storeregister[29][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N1
dffeas \storeregister[25][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][12] .is_wysiwyg = "true";
defparam \storeregister[25][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N11
dffeas \storeregister[17][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][12] .is_wysiwyg = "true";
defparam \storeregister[17][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N11
dffeas \storeregister[21][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][12] .is_wysiwyg = "true";
defparam \storeregister[21][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N10
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[21][12]~q ))) # (!temp_imemload_output_23 & (\storeregister[17][12]~q ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[17][12]~q ),
	.datac(\storeregister[21][12]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hFA44;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N0
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (temp_imemload_output_24 & ((\Mux19~0_combout  & (\storeregister[29][12]~q )) # (!\Mux19~0_combout  & ((\storeregister[25][12]~q ))))) # (!temp_imemload_output_24 & (((\Mux19~0_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[29][12]~q ),
	.datac(\storeregister[25][12]~q ),
	.datad(\Mux19~0_combout ),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hDDA0;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N19
dffeas \storeregister[26][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][12] .is_wysiwyg = "true";
defparam \storeregister[26][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N5
dffeas \storeregister[18][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][12] .is_wysiwyg = "true";
defparam \storeregister[18][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N18
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[26][12]~q )) # (!temp_imemload_output_24 & ((\storeregister[18][12]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[26][12]~q ),
	.datad(\storeregister[18][12]~q ),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hD9C8;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N13
dffeas \storeregister[22][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][12] .is_wysiwyg = "true";
defparam \storeregister[22][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N2
cycloneive_lcell_comb \storeregister[30][12]~feeder (
// Equation(s):
// \storeregister[30][12]~feeder_combout  = Mux19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux19),
	.cin(gnd),
	.combout(\storeregister[30][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][12]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[30][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N3
dffeas \storeregister[30][12] (
	.clk(!CLK),
	.d(\storeregister[30][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][12] .is_wysiwyg = "true";
defparam \storeregister[30][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N12
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = (temp_imemload_output_23 & ((\Mux19~2_combout  & ((\storeregister[30][12]~q ))) # (!\Mux19~2_combout  & (\storeregister[22][12]~q )))) # (!temp_imemload_output_23 & (\Mux19~2_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux19~2_combout ),
	.datac(\storeregister[22][12]~q ),
	.datad(\storeregister[30][12]~q ),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'hEC64;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N15
dffeas \storeregister[16][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][12] .is_wysiwyg = "true";
defparam \storeregister[16][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N28
cycloneive_lcell_comb \storeregister[24][12]~feeder (
// Equation(s):
// \storeregister[24][12]~feeder_combout  = Mux19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux19),
	.cin(gnd),
	.combout(\storeregister[24][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][12]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[24][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N29
dffeas \storeregister[24][12] (
	.clk(!CLK),
	.d(\storeregister[24][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][12] .is_wysiwyg = "true";
defparam \storeregister[24][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N14
cycloneive_lcell_comb \Mux19~4 (
// Equation(s):
// \Mux19~4_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[24][12]~q ))) # (!temp_imemload_output_24 & (\storeregister[16][12]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][12]~q ),
	.datad(\storeregister[24][12]~q ),
	.cin(gnd),
	.combout(\Mux19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~4 .lut_mask = 16'hDC98;
defparam \Mux19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N4
cycloneive_lcell_comb \storeregister[28][12]~feeder (
// Equation(s):
// \storeregister[28][12]~feeder_combout  = Mux19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux19),
	.cin(gnd),
	.combout(\storeregister[28][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][12]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[28][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N5
dffeas \storeregister[28][12] (
	.clk(!CLK),
	.d(\storeregister[28][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][12] .is_wysiwyg = "true";
defparam \storeregister[28][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N29
dffeas \storeregister[20][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][12] .is_wysiwyg = "true";
defparam \storeregister[20][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N30
cycloneive_lcell_comb \Mux19~5 (
// Equation(s):
// \Mux19~5_combout  = (temp_imemload_output_23 & ((\Mux19~4_combout  & (\storeregister[28][12]~q )) # (!\Mux19~4_combout  & ((\storeregister[20][12]~q ))))) # (!temp_imemload_output_23 & (\Mux19~4_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux19~4_combout ),
	.datac(\storeregister[28][12]~q ),
	.datad(\storeregister[20][12]~q ),
	.cin(gnd),
	.combout(\Mux19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~5 .lut_mask = 16'hE6C4;
defparam \Mux19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N8
cycloneive_lcell_comb \Mux19~6 (
// Equation(s):
// \Mux19~6_combout  = (temp_imemload_output_22 & ((\Mux19~3_combout ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((\Mux19~5_combout  & !temp_imemload_output_21))))

	.dataa(temp_imemload_output_22),
	.datab(\Mux19~3_combout ),
	.datac(\Mux19~5_combout ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~6 .lut_mask = 16'hAAD8;
defparam \Mux19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N22
cycloneive_lcell_comb \storeregister[19][12]~feeder (
// Equation(s):
// \storeregister[19][12]~feeder_combout  = Mux19

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux19),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[19][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[19][12]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[19][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N23
dffeas \storeregister[19][12] (
	.clk(!CLK),
	.d(\storeregister[19][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][12] .is_wysiwyg = "true";
defparam \storeregister[19][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N15
dffeas \storeregister[23][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][12] .is_wysiwyg = "true";
defparam \storeregister[23][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N8
cycloneive_lcell_comb \Mux19~7 (
// Equation(s):
// \Mux19~7_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\storeregister[23][12]~q )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & (\storeregister[19][12]~q )))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[19][12]~q ),
	.datad(\storeregister[23][12]~q ),
	.cin(gnd),
	.combout(\Mux19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~7 .lut_mask = 16'hBA98;
defparam \Mux19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N20
cycloneive_lcell_comb \storeregister[31][12]~feeder (
// Equation(s):
// \storeregister[31][12]~feeder_combout  = Mux19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux19),
	.cin(gnd),
	.combout(\storeregister[31][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][12]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[31][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N21
dffeas \storeregister[31][12] (
	.clk(!CLK),
	.d(\storeregister[31][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][12] .is_wysiwyg = "true";
defparam \storeregister[31][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N28
cycloneive_lcell_comb \storeregister[27][12]~feeder (
// Equation(s):
// \storeregister[27][12]~feeder_combout  = Mux19

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux19),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][12]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N29
dffeas \storeregister[27][12] (
	.clk(!CLK),
	.d(\storeregister[27][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][12] .is_wysiwyg = "true";
defparam \storeregister[27][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N2
cycloneive_lcell_comb \Mux19~8 (
// Equation(s):
// \Mux19~8_combout  = (\Mux19~7_combout  & ((\storeregister[31][12]~q ) # ((!temp_imemload_output_24)))) # (!\Mux19~7_combout  & (((temp_imemload_output_24 & \storeregister[27][12]~q ))))

	.dataa(\Mux19~7_combout ),
	.datab(\storeregister[31][12]~q ),
	.datac(temp_imemload_output_24),
	.datad(\storeregister[27][12]~q ),
	.cin(gnd),
	.combout(\Mux19~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~8 .lut_mask = 16'hDA8A;
defparam \Mux19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N19
dffeas \storeregister[7][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][12] .is_wysiwyg = "true";
defparam \storeregister[7][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N21
dffeas \storeregister[6][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][12] .is_wysiwyg = "true";
defparam \storeregister[6][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N18
cycloneive_lcell_comb \Mux19~13 (
// Equation(s):
// \Mux19~13_combout  = (\Mux19~12_combout  & (((\storeregister[7][12]~q )) # (!temp_imemload_output_22))) # (!\Mux19~12_combout  & (temp_imemload_output_22 & ((\storeregister[6][12]~q ))))

	.dataa(\Mux19~12_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[7][12]~q ),
	.datad(\storeregister[6][12]~q ),
	.cin(gnd),
	.combout(\Mux19~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~13 .lut_mask = 16'hE6A2;
defparam \Mux19~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N3
dffeas \storeregister[1][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][12] .is_wysiwyg = "true";
defparam \storeregister[1][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N25
dffeas \storeregister[3][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][12] .is_wysiwyg = "true";
defparam \storeregister[3][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N24
cycloneive_lcell_comb \Mux19~14 (
// Equation(s):
// \Mux19~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][12]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][12]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[1][12]~q ),
	.datac(\storeregister[3][12]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux19~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~14 .lut_mask = 16'hA088;
defparam \Mux19~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N0
cycloneive_lcell_comb \storeregister[2][12]~feeder (
// Equation(s):
// \storeregister[2][12]~feeder_combout  = Mux19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux19),
	.cin(gnd),
	.combout(\storeregister[2][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[2][12]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[2][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N1
dffeas \storeregister[2][12] (
	.clk(!CLK),
	.d(\storeregister[2][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][12] .is_wysiwyg = "true";
defparam \storeregister[2][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N2
cycloneive_lcell_comb \Mux19~15 (
// Equation(s):
// \Mux19~15_combout  = (\Mux19~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][12]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\Mux19~14_combout ),
	.datad(\storeregister[2][12]~q ),
	.cin(gnd),
	.combout(\Mux19~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~15 .lut_mask = 16'hF4F0;
defparam \Mux19~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N6
cycloneive_lcell_comb \Mux19~16 (
// Equation(s):
// \Mux19~16_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\Mux19~13_combout )) # (!temp_imemload_output_23 & ((\Mux19~15_combout )))))

	.dataa(\Mux19~13_combout ),
	.datab(temp_imemload_output_24),
	.datac(temp_imemload_output_23),
	.datad(\Mux19~15_combout ),
	.cin(gnd),
	.combout(\Mux19~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~16 .lut_mask = 16'hE3E0;
defparam \Mux19~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N26
cycloneive_lcell_comb \storeregister[15][12]~feeder (
// Equation(s):
// \storeregister[15][12]~feeder_combout  = Mux19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux19),
	.cin(gnd),
	.combout(\storeregister[15][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][12]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N27
dffeas \storeregister[15][12] (
	.clk(!CLK),
	.d(\storeregister[15][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][12] .is_wysiwyg = "true";
defparam \storeregister[15][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N0
cycloneive_lcell_comb \storeregister[14][12]~feeder (
// Equation(s):
// \storeregister[14][12]~feeder_combout  = Mux19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux19),
	.cin(gnd),
	.combout(\storeregister[14][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][12]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N1
dffeas \storeregister[14][12] (
	.clk(!CLK),
	.d(\storeregister[14][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][12] .is_wysiwyg = "true";
defparam \storeregister[14][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N11
dffeas \storeregister[13][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][12] .is_wysiwyg = "true";
defparam \storeregister[13][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N25
dffeas \storeregister[12][12] (
	.clk(!CLK),
	.d(Mux19),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][12] .is_wysiwyg = "true";
defparam \storeregister[12][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N10
cycloneive_lcell_comb \Mux19~17 (
// Equation(s):
// \Mux19~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][12]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[12][12]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[13][12]~q ),
	.datad(\storeregister[12][12]~q ),
	.cin(gnd),
	.combout(\Mux19~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~17 .lut_mask = 16'hB9A8;
defparam \Mux19~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N8
cycloneive_lcell_comb \Mux19~18 (
// Equation(s):
// \Mux19~18_combout  = (temp_imemload_output_22 & ((\Mux19~17_combout  & (\storeregister[15][12]~q )) # (!\Mux19~17_combout  & ((\storeregister[14][12]~q ))))) # (!temp_imemload_output_22 & (((\Mux19~17_combout ))))

	.dataa(\storeregister[15][12]~q ),
	.datab(\storeregister[14][12]~q ),
	.datac(temp_imemload_output_22),
	.datad(\Mux19~17_combout ),
	.cin(gnd),
	.combout(\Mux19~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~18 .lut_mask = 16'hAFC0;
defparam \Mux19~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N11
dffeas \storeregister[10][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][12] .is_wysiwyg = "true";
defparam \storeregister[10][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N25
dffeas \storeregister[8][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][12] .is_wysiwyg = "true";
defparam \storeregister[8][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N10
cycloneive_lcell_comb \Mux19~10 (
// Equation(s):
// \Mux19~10_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\storeregister[10][12]~q )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & ((\storeregister[8][12]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[10][12]~q ),
	.datad(\storeregister[8][12]~q ),
	.cin(gnd),
	.combout(\Mux19~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~10 .lut_mask = 16'hB9A8;
defparam \Mux19~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N23
dffeas \storeregister[9][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][12] .is_wysiwyg = "true";
defparam \storeregister[9][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N21
dffeas \storeregister[11][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][12] .is_wysiwyg = "true";
defparam \storeregister[11][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N22
cycloneive_lcell_comb \Mux19~11 (
// Equation(s):
// \Mux19~11_combout  = (\Mux19~10_combout  & (((\storeregister[11][12]~q )) # (!temp_imemload_output_21))) # (!\Mux19~10_combout  & (temp_imemload_output_21 & (\storeregister[9][12]~q )))

	.dataa(\Mux19~10_combout ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[9][12]~q ),
	.datad(\storeregister[11][12]~q ),
	.cin(gnd),
	.combout(\Mux19~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~11 .lut_mask = 16'hEA62;
defparam \Mux19~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N3
dffeas \storeregister[28][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][10] .is_wysiwyg = "true";
defparam \storeregister[28][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N25
dffeas \storeregister[20][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][10] .is_wysiwyg = "true";
defparam \storeregister[20][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N2
cycloneive_lcell_comb \Mux21~5 (
// Equation(s):
// \Mux21~5_combout  = (\Mux21~4_combout  & (((\storeregister[28][10]~q )) # (!temp_imemload_output_23))) # (!\Mux21~4_combout  & (temp_imemload_output_23 & ((\storeregister[20][10]~q ))))

	.dataa(\Mux21~4_combout ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[28][10]~q ),
	.datad(\storeregister[20][10]~q ),
	.cin(gnd),
	.combout(\Mux21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~5 .lut_mask = 16'hE6A2;
defparam \Mux21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N25
dffeas \storeregister[26][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][10] .is_wysiwyg = "true";
defparam \storeregister[26][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N24
cycloneive_lcell_comb \Mux21~2 (
// Equation(s):
// \Mux21~2_combout  = (temp_imemload_output_24 & (((\storeregister[26][10]~q ) # (temp_imemload_output_23)))) # (!temp_imemload_output_24 & (\storeregister[18][10]~q  & ((!temp_imemload_output_23))))

	.dataa(\storeregister[18][10]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[26][10]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~2 .lut_mask = 16'hCCE2;
defparam \Mux21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N27
dffeas \storeregister[22][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][10] .is_wysiwyg = "true";
defparam \storeregister[22][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N1
dffeas \storeregister[30][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][10] .is_wysiwyg = "true";
defparam \storeregister[30][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N26
cycloneive_lcell_comb \Mux21~3 (
// Equation(s):
// \Mux21~3_combout  = (temp_imemload_output_23 & ((\Mux21~2_combout  & ((\storeregister[30][10]~q ))) # (!\Mux21~2_combout  & (\storeregister[22][10]~q )))) # (!temp_imemload_output_23 & (\Mux21~2_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux21~2_combout ),
	.datac(\storeregister[22][10]~q ),
	.datad(\storeregister[30][10]~q ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~3 .lut_mask = 16'hEC64;
defparam \Mux21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N0
cycloneive_lcell_comb \Mux21~6 (
// Equation(s):
// \Mux21~6_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22)))) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & ((\Mux21~3_combout ))) # (!temp_imemload_output_22 & (\Mux21~5_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux21~5_combout ),
	.datac(temp_imemload_output_22),
	.datad(\Mux21~3_combout ),
	.cin(gnd),
	.combout(\Mux21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~6 .lut_mask = 16'hF4A4;
defparam \Mux21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N12
cycloneive_lcell_comb \storeregister[21][10]~feeder (
// Equation(s):
// \storeregister[21][10]~feeder_combout  = Mux21

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux21),
	.cin(gnd),
	.combout(\storeregister[21][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][10]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[21][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N13
dffeas \storeregister[21][10] (
	.clk(!CLK),
	.d(\storeregister[21][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][10] .is_wysiwyg = "true";
defparam \storeregister[21][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N27
dffeas \storeregister[17][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][10] .is_wysiwyg = "true";
defparam \storeregister[17][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N26
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (temp_imemload_output_23 & ((\storeregister[21][10]~q ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\storeregister[17][10]~q  & !temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[21][10]~q ),
	.datac(\storeregister[17][10]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hAAD8;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N11
dffeas \storeregister[25][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][10] .is_wysiwyg = "true";
defparam \storeregister[25][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N25
dffeas \storeregister[29][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][10] .is_wysiwyg = "true";
defparam \storeregister[29][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N10
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (temp_imemload_output_24 & ((\Mux21~0_combout  & ((\storeregister[29][10]~q ))) # (!\Mux21~0_combout  & (\storeregister[25][10]~q )))) # (!temp_imemload_output_24 & (\Mux21~0_combout ))

	.dataa(temp_imemload_output_24),
	.datab(\Mux21~0_combout ),
	.datac(\storeregister[25][10]~q ),
	.datad(\storeregister[29][10]~q ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hEC64;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N15
dffeas \storeregister[19][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][10] .is_wysiwyg = "true";
defparam \storeregister[19][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N13
dffeas \storeregister[23][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][10] .is_wysiwyg = "true";
defparam \storeregister[23][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N14
cycloneive_lcell_comb \Mux21~7 (
// Equation(s):
// \Mux21~7_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[23][10]~q ))) # (!temp_imemload_output_23 & (\storeregister[19][10]~q ))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[19][10]~q ),
	.datad(\storeregister[23][10]~q ),
	.cin(gnd),
	.combout(\Mux21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~7 .lut_mask = 16'hDC98;
defparam \Mux21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N5
dffeas \storeregister[27][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][10] .is_wysiwyg = "true";
defparam \storeregister[27][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N8
cycloneive_lcell_comb \storeregister[31][10]~feeder (
// Equation(s):
// \storeregister[31][10]~feeder_combout  = Mux21

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux21),
	.cin(gnd),
	.combout(\storeregister[31][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][10]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[31][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N9
dffeas \storeregister[31][10] (
	.clk(!CLK),
	.d(\storeregister[31][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][10] .is_wysiwyg = "true";
defparam \storeregister[31][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N4
cycloneive_lcell_comb \Mux21~8 (
// Equation(s):
// \Mux21~8_combout  = (\Mux21~7_combout  & (((\storeregister[31][10]~q )) # (!temp_imemload_output_24))) # (!\Mux21~7_combout  & (temp_imemload_output_24 & (\storeregister[27][10]~q )))

	.dataa(\Mux21~7_combout ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[27][10]~q ),
	.datad(\storeregister[31][10]~q ),
	.cin(gnd),
	.combout(\Mux21~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~8 .lut_mask = 16'hEA62;
defparam \Mux21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N12
cycloneive_lcell_comb \storeregister[8][10]~feeder (
// Equation(s):
// \storeregister[8][10]~feeder_combout  = Mux21

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux21),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[8][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[8][10]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[8][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N13
dffeas \storeregister[8][10] (
	.clk(!CLK),
	.d(\storeregister[8][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][10] .is_wysiwyg = "true";
defparam \storeregister[8][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y39_N25
dffeas \storeregister[10][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][10] .is_wysiwyg = "true";
defparam \storeregister[10][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N26
cycloneive_lcell_comb \Mux21~10 (
// Equation(s):
// \Mux21~10_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[10][10]~q ))) # (!temp_imemload_output_22 & (\storeregister[8][10]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[8][10]~q ),
	.datad(\storeregister[10][10]~q ),
	.cin(gnd),
	.combout(\Mux21~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~10 .lut_mask = 16'hDC98;
defparam \Mux21~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N15
dffeas \storeregister[9][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][10] .is_wysiwyg = "true";
defparam \storeregister[9][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N1
dffeas \storeregister[11][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][10] .is_wysiwyg = "true";
defparam \storeregister[11][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N14
cycloneive_lcell_comb \Mux21~11 (
// Equation(s):
// \Mux21~11_combout  = (temp_imemload_output_21 & ((\Mux21~10_combout  & ((\storeregister[11][10]~q ))) # (!\Mux21~10_combout  & (\storeregister[9][10]~q )))) # (!temp_imemload_output_21 & (\Mux21~10_combout ))

	.dataa(temp_imemload_output_21),
	.datab(\Mux21~10_combout ),
	.datac(\storeregister[9][10]~q ),
	.datad(\storeregister[11][10]~q ),
	.cin(gnd),
	.combout(\Mux21~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~11 .lut_mask = 16'hEC64;
defparam \Mux21~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N31
dffeas \storeregister[7][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][10] .is_wysiwyg = "true";
defparam \storeregister[7][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y41_N19
dffeas \storeregister[4][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][10] .is_wysiwyg = "true";
defparam \storeregister[4][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y41_N9
dffeas \storeregister[5][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][10] .is_wysiwyg = "true";
defparam \storeregister[5][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N8
cycloneive_lcell_comb \Mux21~12 (
// Equation(s):
// \Mux21~12_combout  = (temp_imemload_output_21 & (((\storeregister[5][10]~q ) # (temp_imemload_output_22)))) # (!temp_imemload_output_21 & (\storeregister[4][10]~q  & ((!temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[4][10]~q ),
	.datac(\storeregister[5][10]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux21~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~12 .lut_mask = 16'hAAE4;
defparam \Mux21~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N30
cycloneive_lcell_comb \Mux21~13 (
// Equation(s):
// \Mux21~13_combout  = (temp_imemload_output_22 & ((\Mux21~12_combout  & ((\storeregister[7][10]~q ))) # (!\Mux21~12_combout  & (\storeregister[6][10]~q )))) # (!temp_imemload_output_22 & (((\Mux21~12_combout ))))

	.dataa(\storeregister[6][10]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[7][10]~q ),
	.datad(\Mux21~12_combout ),
	.cin(gnd),
	.combout(\Mux21~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~13 .lut_mask = 16'hF388;
defparam \Mux21~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N20
cycloneive_lcell_comb \storeregister[2][10]~feeder (
// Equation(s):
// \storeregister[2][10]~feeder_combout  = Mux21

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux21),
	.cin(gnd),
	.combout(\storeregister[2][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[2][10]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[2][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N21
dffeas \storeregister[2][10] (
	.clk(!CLK),
	.d(\storeregister[2][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][10] .is_wysiwyg = "true";
defparam \storeregister[2][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N25
dffeas \storeregister[3][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][10] .is_wysiwyg = "true";
defparam \storeregister[3][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N24
cycloneive_lcell_comb \Mux21~14 (
// Equation(s):
// \Mux21~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][10]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][10]~q ))))

	.dataa(\storeregister[1][10]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[3][10]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux21~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~14 .lut_mask = 16'hE200;
defparam \Mux21~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N26
cycloneive_lcell_comb \Mux21~15 (
// Equation(s):
// \Mux21~15_combout  = (\Mux21~14_combout ) # ((!temp_imemload_output_21 & (\storeregister[2][10]~q  & temp_imemload_output_22)))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[2][10]~q ),
	.datac(\Mux21~14_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux21~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~15 .lut_mask = 16'hF4F0;
defparam \Mux21~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N22
cycloneive_lcell_comb \Mux21~16 (
// Equation(s):
// \Mux21~16_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\Mux21~13_combout )) # (!temp_imemload_output_23 & ((\Mux21~15_combout )))))

	.dataa(\Mux21~13_combout ),
	.datab(temp_imemload_output_24),
	.datac(temp_imemload_output_23),
	.datad(\Mux21~15_combout ),
	.cin(gnd),
	.combout(\Mux21~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~16 .lut_mask = 16'hE3E0;
defparam \Mux21~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N27
dffeas \storeregister[12][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][10] .is_wysiwyg = "true";
defparam \storeregister[12][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N13
dffeas \storeregister[13][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][10] .is_wysiwyg = "true";
defparam \storeregister[13][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N26
cycloneive_lcell_comb \Mux21~17 (
// Equation(s):
// \Mux21~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][10]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[12][10]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[12][10]~q ),
	.datad(\storeregister[13][10]~q ),
	.cin(gnd),
	.combout(\Mux21~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~17 .lut_mask = 16'hBA98;
defparam \Mux21~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N16
cycloneive_lcell_comb \storeregister[14][10]~feeder (
// Equation(s):
// \storeregister[14][10]~feeder_combout  = Mux21

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux21),
	.cin(gnd),
	.combout(\storeregister[14][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][10]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N17
dffeas \storeregister[14][10] (
	.clk(!CLK),
	.d(\storeregister[14][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][10] .is_wysiwyg = "true";
defparam \storeregister[14][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N29
dffeas \storeregister[15][10] (
	.clk(!CLK),
	.d(Mux21),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][10] .is_wysiwyg = "true";
defparam \storeregister[15][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N12
cycloneive_lcell_comb \Mux21~18 (
// Equation(s):
// \Mux21~18_combout  = (\Mux21~17_combout  & (((\storeregister[15][10]~q ) # (!temp_imemload_output_22)))) # (!\Mux21~17_combout  & (\storeregister[14][10]~q  & (temp_imemload_output_22)))

	.dataa(\Mux21~17_combout ),
	.datab(\storeregister[14][10]~q ),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[15][10]~q ),
	.cin(gnd),
	.combout(\Mux21~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~18 .lut_mask = 16'hEA4A;
defparam \Mux21~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N9
dffeas \storeregister[26][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][11] .is_wysiwyg = "true";
defparam \storeregister[26][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N1
dffeas \storeregister[22][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][11] .is_wysiwyg = "true";
defparam \storeregister[22][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N19
dffeas \storeregister[18][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][11] .is_wysiwyg = "true";
defparam \storeregister[18][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N18
cycloneive_lcell_comb \Mux20~2 (
// Equation(s):
// \Mux20~2_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[22][11]~q )) # (!temp_imemload_output_23 & ((\storeregister[18][11]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[22][11]~q ),
	.datac(\storeregister[18][11]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~2 .lut_mask = 16'hEE50;
defparam \Mux20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N26
cycloneive_lcell_comb \Mux20~3 (
// Equation(s):
// \Mux20~3_combout  = (temp_imemload_output_24 & ((\Mux20~2_combout  & (\storeregister[30][11]~q )) # (!\Mux20~2_combout  & ((\storeregister[26][11]~q ))))) # (!temp_imemload_output_24 & (((\Mux20~2_combout ))))

	.dataa(\storeregister[30][11]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[26][11]~q ),
	.datad(\Mux20~2_combout ),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~3 .lut_mask = 16'hBBC0;
defparam \Mux20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N22
cycloneive_lcell_comb \storeregister[28][11]~feeder (
// Equation(s):
// \storeregister[28][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux20),
	.cin(gnd),
	.combout(\storeregister[28][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][11]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[28][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N23
dffeas \storeregister[28][11] (
	.clk(!CLK),
	.d(\storeregister[28][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][11] .is_wysiwyg = "true";
defparam \storeregister[28][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N21
dffeas \storeregister[16][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][11] .is_wysiwyg = "true";
defparam \storeregister[16][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N20
cycloneive_lcell_comb \Mux20~4 (
// Equation(s):
// \Mux20~4_combout  = (temp_imemload_output_23 & ((\storeregister[20][11]~q ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\storeregister[16][11]~q  & !temp_imemload_output_24))))

	.dataa(\storeregister[20][11]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[16][11]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~4 .lut_mask = 16'hCCB8;
defparam \Mux20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N0
cycloneive_lcell_comb \Mux20~5 (
// Equation(s):
// \Mux20~5_combout  = (temp_imemload_output_24 & ((\Mux20~4_combout  & ((\storeregister[28][11]~q ))) # (!\Mux20~4_combout  & (\storeregister[24][11]~q )))) # (!temp_imemload_output_24 & (((\Mux20~4_combout ))))

	.dataa(\storeregister[24][11]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[28][11]~q ),
	.datad(\Mux20~4_combout ),
	.cin(gnd),
	.combout(\Mux20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~5 .lut_mask = 16'hF388;
defparam \Mux20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N10
cycloneive_lcell_comb \Mux20~6 (
// Equation(s):
// \Mux20~6_combout  = (temp_imemload_output_22 & ((\Mux20~3_combout ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((\Mux20~5_combout  & !temp_imemload_output_21))))

	.dataa(\Mux20~3_combout ),
	.datab(\Mux20~5_combout ),
	.datac(temp_imemload_output_22),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~6 .lut_mask = 16'hF0AC;
defparam \Mux20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N4
cycloneive_lcell_comb \storeregister[21][11]~feeder (
// Equation(s):
// \storeregister[21][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux20),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[21][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][11]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[21][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N5
dffeas \storeregister[21][11] (
	.clk(!CLK),
	.d(\storeregister[21][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][11] .is_wysiwyg = "true";
defparam \storeregister[21][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N14
cycloneive_lcell_comb \storeregister[29][11]~feeder (
// Equation(s):
// \storeregister[29][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux20),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[29][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][11]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[29][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N15
dffeas \storeregister[29][11] (
	.clk(!CLK),
	.d(\storeregister[29][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][11] .is_wysiwyg = "true";
defparam \storeregister[29][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N17
dffeas \storeregister[25][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][11] .is_wysiwyg = "true";
defparam \storeregister[25][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N24
cycloneive_lcell_comb \storeregister[17][11]~feeder (
// Equation(s):
// \storeregister[17][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux20),
	.cin(gnd),
	.combout(\storeregister[17][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[17][11]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[17][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N25
dffeas \storeregister[17][11] (
	.clk(!CLK),
	.d(\storeregister[17][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][11] .is_wysiwyg = "true";
defparam \storeregister[17][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N16
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (temp_imemload_output_24 & ((temp_imemload_output_23) # ((\storeregister[25][11]~q )))) # (!temp_imemload_output_24 & (!temp_imemload_output_23 & ((\storeregister[17][11]~q ))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[25][11]~q ),
	.datad(\storeregister[17][11]~q ),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hB9A8;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N10
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (temp_imemload_output_23 & ((\Mux20~0_combout  & ((\storeregister[29][11]~q ))) # (!\Mux20~0_combout  & (\storeregister[21][11]~q )))) # (!temp_imemload_output_23 & (((\Mux20~0_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[21][11]~q ),
	.datac(\storeregister[29][11]~q ),
	.datad(\Mux20~0_combout ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hF588;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N28
cycloneive_lcell_comb \storeregister[31][11]~feeder (
// Equation(s):
// \storeregister[31][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux20),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[31][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][11]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[31][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N29
dffeas \storeregister[31][11] (
	.clk(!CLK),
	.d(\storeregister[31][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][11] .is_wysiwyg = "true";
defparam \storeregister[31][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N2
cycloneive_lcell_comb \storeregister[19][11]~feeder (
// Equation(s):
// \storeregister[19][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux20),
	.cin(gnd),
	.combout(\storeregister[19][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[19][11]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[19][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N3
dffeas \storeregister[19][11] (
	.clk(!CLK),
	.d(\storeregister[19][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][11] .is_wysiwyg = "true";
defparam \storeregister[19][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N26
cycloneive_lcell_comb \Mux20~7 (
// Equation(s):
// \Mux20~7_combout  = (temp_imemload_output_24 & ((\storeregister[27][11]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[19][11]~q  & !temp_imemload_output_23))))

	.dataa(\storeregister[27][11]~q ),
	.datab(\storeregister[19][11]~q ),
	.datac(temp_imemload_output_24),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~7 .lut_mask = 16'hF0AC;
defparam \Mux20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N3
dffeas \storeregister[23][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][11] .is_wysiwyg = "true";
defparam \storeregister[23][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N18
cycloneive_lcell_comb \Mux20~8 (
// Equation(s):
// \Mux20~8_combout  = (temp_imemload_output_23 & ((\Mux20~7_combout  & (\storeregister[31][11]~q )) # (!\Mux20~7_combout  & ((\storeregister[23][11]~q ))))) # (!temp_imemload_output_23 & (((\Mux20~7_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[31][11]~q ),
	.datac(\Mux20~7_combout ),
	.datad(\storeregister[23][11]~q ),
	.cin(gnd),
	.combout(\Mux20~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~8 .lut_mask = 16'hDAD0;
defparam \Mux20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N8
cycloneive_lcell_comb \storeregister[7][11]~feeder (
// Equation(s):
// \storeregister[7][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux20),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[7][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[7][11]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[7][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N9
dffeas \storeregister[7][11] (
	.clk(!CLK),
	.d(\storeregister[7][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][11] .is_wysiwyg = "true";
defparam \storeregister[7][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y42_N9
dffeas \storeregister[5][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][11] .is_wysiwyg = "true";
defparam \storeregister[5][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y42_N7
dffeas \storeregister[4][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][11] .is_wysiwyg = "true";
defparam \storeregister[4][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N8
cycloneive_lcell_comb \Mux20~10 (
// Equation(s):
// \Mux20~10_combout  = (temp_imemload_output_22 & (temp_imemload_output_21)) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & (\storeregister[5][11]~q )) # (!temp_imemload_output_21 & ((\storeregister[4][11]~q )))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[5][11]~q ),
	.datad(\storeregister[4][11]~q ),
	.cin(gnd),
	.combout(\Mux20~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~10 .lut_mask = 16'hD9C8;
defparam \Mux20~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N4
cycloneive_lcell_comb \storeregister[6][11]~feeder (
// Equation(s):
// \storeregister[6][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux20),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[6][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[6][11]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[6][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N5
dffeas \storeregister[6][11] (
	.clk(!CLK),
	.d(\storeregister[6][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][11] .is_wysiwyg = "true";
defparam \storeregister[6][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N6
cycloneive_lcell_comb \Mux20~11 (
// Equation(s):
// \Mux20~11_combout  = (\Mux20~10_combout  & ((\storeregister[7][11]~q ) # ((!temp_imemload_output_22)))) # (!\Mux20~10_combout  & (((\storeregister[6][11]~q  & temp_imemload_output_22))))

	.dataa(\storeregister[7][11]~q ),
	.datab(\Mux20~10_combout ),
	.datac(\storeregister[6][11]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux20~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~11 .lut_mask = 16'hB8CC;
defparam \Mux20~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N1
dffeas \storeregister[3][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][11] .is_wysiwyg = "true";
defparam \storeregister[3][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N0
cycloneive_lcell_comb \Mux20~14 (
// Equation(s):
// \Mux20~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][11]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][11]~q ))))

	.dataa(\storeregister[1][11]~q ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[3][11]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux20~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~14 .lut_mask = 16'hC088;
defparam \Mux20~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N5
dffeas \storeregister[2][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][11] .is_wysiwyg = "true";
defparam \storeregister[2][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N4
cycloneive_lcell_comb \Mux20~15 (
// Equation(s):
// \Mux20~15_combout  = (\Mux20~14_combout ) # ((!temp_imemload_output_21 & (\storeregister[2][11]~q  & temp_imemload_output_22)))

	.dataa(temp_imemload_output_21),
	.datab(\Mux20~14_combout ),
	.datac(\storeregister[2][11]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux20~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~15 .lut_mask = 16'hDCCC;
defparam \Mux20~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N4
cycloneive_lcell_comb \storeregister[11][11]~feeder (
// Equation(s):
// \storeregister[11][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux20),
	.cin(gnd),
	.combout(\storeregister[11][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[11][11]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[11][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N5
dffeas \storeregister[11][11] (
	.clk(!CLK),
	.d(\storeregister[11][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][11] .is_wysiwyg = "true";
defparam \storeregister[11][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N14
cycloneive_lcell_comb \storeregister[9][11]~feeder (
// Equation(s):
// \storeregister[9][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux20),
	.cin(gnd),
	.combout(\storeregister[9][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[9][11]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[9][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N15
dffeas \storeregister[9][11] (
	.clk(!CLK),
	.d(\storeregister[9][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][11] .is_wysiwyg = "true";
defparam \storeregister[9][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N30
cycloneive_lcell_comb \Mux20~13 (
// Equation(s):
// \Mux20~13_combout  = (\Mux20~12_combout  & ((\storeregister[11][11]~q ) # ((!temp_imemload_output_21)))) # (!\Mux20~12_combout  & (((\storeregister[9][11]~q  & temp_imemload_output_21))))

	.dataa(\Mux20~12_combout ),
	.datab(\storeregister[11][11]~q ),
	.datac(\storeregister[9][11]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux20~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~13 .lut_mask = 16'hD8AA;
defparam \Mux20~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N24
cycloneive_lcell_comb \Mux20~16 (
// Equation(s):
// \Mux20~16_combout  = (temp_imemload_output_24 & ((temp_imemload_output_23) # ((\Mux20~13_combout )))) # (!temp_imemload_output_24 & (!temp_imemload_output_23 & (\Mux20~15_combout )))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\Mux20~15_combout ),
	.datad(\Mux20~13_combout ),
	.cin(gnd),
	.combout(\Mux20~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~16 .lut_mask = 16'hBA98;
defparam \Mux20~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N18
cycloneive_lcell_comb \storeregister[15][11]~feeder (
// Equation(s):
// \storeregister[15][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux20),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[15][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][11]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[15][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N19
dffeas \storeregister[15][11] (
	.clk(!CLK),
	.d(\storeregister[15][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][11] .is_wysiwyg = "true";
defparam \storeregister[15][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N14
cycloneive_lcell_comb \storeregister[14][11]~feeder (
// Equation(s):
// \storeregister[14][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux20),
	.cin(gnd),
	.combout(\storeregister[14][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][11]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N15
dffeas \storeregister[14][11] (
	.clk(!CLK),
	.d(\storeregister[14][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][11] .is_wysiwyg = "true";
defparam \storeregister[14][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N9
dffeas \storeregister[13][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][11] .is_wysiwyg = "true";
defparam \storeregister[13][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N7
dffeas \storeregister[12][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][11] .is_wysiwyg = "true";
defparam \storeregister[12][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N6
cycloneive_lcell_comb \Mux20~17 (
// Equation(s):
// \Mux20~17_combout  = (temp_imemload_output_21 & ((\storeregister[13][11]~q ) # ((temp_imemload_output_22)))) # (!temp_imemload_output_21 & (((\storeregister[12][11]~q  & !temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[13][11]~q ),
	.datac(\storeregister[12][11]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux20~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~17 .lut_mask = 16'hAAD8;
defparam \Mux20~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N2
cycloneive_lcell_comb \Mux20~18 (
// Equation(s):
// \Mux20~18_combout  = (\Mux20~17_combout  & ((\storeregister[15][11]~q ) # ((!temp_imemload_output_22)))) # (!\Mux20~17_combout  & (((\storeregister[14][11]~q  & temp_imemload_output_22))))

	.dataa(\storeregister[15][11]~q ),
	.datab(\storeregister[14][11]~q ),
	.datac(\Mux20~17_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux20~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~18 .lut_mask = 16'hACF0;
defparam \Mux20~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N15
dffeas \storeregister[17][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][9] .is_wysiwyg = "true";
defparam \storeregister[17][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N14
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[25][9]~q )) # (!temp_imemload_output_24 & ((\storeregister[17][9]~q )))))

	.dataa(\storeregister[25][9]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[17][9]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hEE30;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N26
cycloneive_lcell_comb \storeregister[29][9]~feeder (
// Equation(s):
// \storeregister[29][9]~feeder_combout  = Mux22

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux22),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[29][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][9]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[29][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N27
dffeas \storeregister[29][9] (
	.clk(!CLK),
	.d(\storeregister[29][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][9] .is_wysiwyg = "true";
defparam \storeregister[29][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N8
cycloneive_lcell_comb \storeregister[21][9]~feeder (
// Equation(s):
// \storeregister[21][9]~feeder_combout  = Mux22

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux22),
	.cin(gnd),
	.combout(\storeregister[21][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][9]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[21][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N9
dffeas \storeregister[21][9] (
	.clk(!CLK),
	.d(\storeregister[21][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][9] .is_wysiwyg = "true";
defparam \storeregister[21][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N0
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (temp_imemload_output_23 & ((\Mux22~0_combout  & (\storeregister[29][9]~q )) # (!\Mux22~0_combout  & ((\storeregister[21][9]~q ))))) # (!temp_imemload_output_23 & (\Mux22~0_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux22~0_combout ),
	.datac(\storeregister[29][9]~q ),
	.datad(\storeregister[21][9]~q ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hE6C4;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N15
dffeas \storeregister[30][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][9] .is_wysiwyg = "true";
defparam \storeregister[30][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N21
dffeas \storeregister[26][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][9] .is_wysiwyg = "true";
defparam \storeregister[26][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N20
cycloneive_lcell_comb \Mux22~3 (
// Equation(s):
// \Mux22~3_combout  = (\Mux22~2_combout  & ((\storeregister[30][9]~q ) # ((!temp_imemload_output_24)))) # (!\Mux22~2_combout  & (((\storeregister[26][9]~q  & temp_imemload_output_24))))

	.dataa(\Mux22~2_combout ),
	.datab(\storeregister[30][9]~q ),
	.datac(\storeregister[26][9]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~3 .lut_mask = 16'hD8AA;
defparam \Mux22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N17
dffeas \storeregister[28][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][9] .is_wysiwyg = "true";
defparam \storeregister[28][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N26
cycloneive_lcell_comb \storeregister[24][9]~feeder (
// Equation(s):
// \storeregister[24][9]~feeder_combout  = Mux22

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux22),
	.cin(gnd),
	.combout(\storeregister[24][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][9]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[24][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N27
dffeas \storeregister[24][9] (
	.clk(!CLK),
	.d(\storeregister[24][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][9] .is_wysiwyg = "true";
defparam \storeregister[24][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N16
cycloneive_lcell_comb \Mux22~5 (
// Equation(s):
// \Mux22~5_combout  = (\Mux22~4_combout  & (((\storeregister[28][9]~q )) # (!temp_imemload_output_24))) # (!\Mux22~4_combout  & (temp_imemload_output_24 & ((\storeregister[24][9]~q ))))

	.dataa(\Mux22~4_combout ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[28][9]~q ),
	.datad(\storeregister[24][9]~q ),
	.cin(gnd),
	.combout(\Mux22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~5 .lut_mask = 16'hE6A2;
defparam \Mux22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N30
cycloneive_lcell_comb \Mux22~6 (
// Equation(s):
// \Mux22~6_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22)))) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\Mux22~3_combout )) # (!temp_imemload_output_22 & ((\Mux22~5_combout )))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux22~3_combout ),
	.datac(temp_imemload_output_22),
	.datad(\Mux22~5_combout ),
	.cin(gnd),
	.combout(\Mux22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~6 .lut_mask = 16'hE5E0;
defparam \Mux22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N9
dffeas \storeregister[23][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][9] .is_wysiwyg = "true";
defparam \storeregister[23][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N25
dffeas \storeregister[31][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][9] .is_wysiwyg = "true";
defparam \storeregister[31][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N27
dffeas \storeregister[19][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][9] .is_wysiwyg = "true";
defparam \storeregister[19][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N30
cycloneive_lcell_comb \storeregister[27][9]~feeder (
// Equation(s):
// \storeregister[27][9]~feeder_combout  = Mux22

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux22),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][9]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N31
dffeas \storeregister[27][9] (
	.clk(!CLK),
	.d(\storeregister[27][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][9] .is_wysiwyg = "true";
defparam \storeregister[27][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N26
cycloneive_lcell_comb \Mux22~7 (
// Equation(s):
// \Mux22~7_combout  = (temp_imemload_output_24 & ((temp_imemload_output_23) # ((\storeregister[27][9]~q )))) # (!temp_imemload_output_24 & (!temp_imemload_output_23 & (\storeregister[19][9]~q )))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[19][9]~q ),
	.datad(\storeregister[27][9]~q ),
	.cin(gnd),
	.combout(\Mux22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~7 .lut_mask = 16'hBA98;
defparam \Mux22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N24
cycloneive_lcell_comb \Mux22~8 (
// Equation(s):
// \Mux22~8_combout  = (temp_imemload_output_23 & ((\Mux22~7_combout  & ((\storeregister[31][9]~q ))) # (!\Mux22~7_combout  & (\storeregister[23][9]~q )))) # (!temp_imemload_output_23 & (((\Mux22~7_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[23][9]~q ),
	.datac(\storeregister[31][9]~q ),
	.datad(\Mux22~7_combout ),
	.cin(gnd),
	.combout(\Mux22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~8 .lut_mask = 16'hF588;
defparam \Mux22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y41_N21
dffeas \storeregister[5][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][9] .is_wysiwyg = "true";
defparam \storeregister[5][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N20
cycloneive_lcell_comb \Mux22~10 (
// Equation(s):
// \Mux22~10_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[5][9]~q ))) # (!temp_imemload_output_21 & (\storeregister[4][9]~q ))))

	.dataa(\storeregister[4][9]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[5][9]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux22~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~10 .lut_mask = 16'hFC22;
defparam \Mux22~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N29
dffeas \storeregister[7][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][9] .is_wysiwyg = "true";
defparam \storeregister[7][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N15
dffeas \storeregister[6][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][9] .is_wysiwyg = "true";
defparam \storeregister[6][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N14
cycloneive_lcell_comb \Mux22~11 (
// Equation(s):
// \Mux22~11_combout  = (\Mux22~10_combout  & ((\storeregister[7][9]~q ) # ((!temp_imemload_output_22)))) # (!\Mux22~10_combout  & (((\storeregister[6][9]~q  & temp_imemload_output_22))))

	.dataa(\Mux22~10_combout ),
	.datab(\storeregister[7][9]~q ),
	.datac(\storeregister[6][9]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux22~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~11 .lut_mask = 16'hD8AA;
defparam \Mux22~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y42_N11
dffeas \storeregister[12][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][9] .is_wysiwyg = "true";
defparam \storeregister[12][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N29
dffeas \storeregister[13][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][9] .is_wysiwyg = "true";
defparam \storeregister[13][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N10
cycloneive_lcell_comb \Mux22~17 (
// Equation(s):
// \Mux22~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][9]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[12][9]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[12][9]~q ),
	.datad(\storeregister[13][9]~q ),
	.cin(gnd),
	.combout(\Mux22~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~17 .lut_mask = 16'hBA98;
defparam \Mux22~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N3
dffeas \storeregister[14][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][9] .is_wysiwyg = "true";
defparam \storeregister[14][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N12
cycloneive_lcell_comb \storeregister[15][9]~feeder (
// Equation(s):
// \storeregister[15][9]~feeder_combout  = Mux22

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux22),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[15][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][9]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[15][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N13
dffeas \storeregister[15][9] (
	.clk(!CLK),
	.d(\storeregister[15][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][9] .is_wysiwyg = "true";
defparam \storeregister[15][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N14
cycloneive_lcell_comb \Mux22~18 (
// Equation(s):
// \Mux22~18_combout  = (\Mux22~17_combout  & (((\storeregister[15][9]~q ) # (!temp_imemload_output_22)))) # (!\Mux22~17_combout  & (\storeregister[14][9]~q  & (temp_imemload_output_22)))

	.dataa(\Mux22~17_combout ),
	.datab(\storeregister[14][9]~q ),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[15][9]~q ),
	.cin(gnd),
	.combout(\Mux22~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~18 .lut_mask = 16'hEA4A;
defparam \Mux22~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N3
dffeas \storeregister[8][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][9] .is_wysiwyg = "true";
defparam \storeregister[8][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N13
dffeas \storeregister[10][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][9] .is_wysiwyg = "true";
defparam \storeregister[10][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N2
cycloneive_lcell_comb \Mux22~12 (
// Equation(s):
// \Mux22~12_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\storeregister[10][9]~q )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & (\storeregister[8][9]~q )))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[8][9]~q ),
	.datad(\storeregister[10][9]~q ),
	.cin(gnd),
	.combout(\Mux22~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~12 .lut_mask = 16'hBA98;
defparam \Mux22~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N13
dffeas \storeregister[11][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][9] .is_wysiwyg = "true";
defparam \storeregister[11][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N3
dffeas \storeregister[9][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][9] .is_wysiwyg = "true";
defparam \storeregister[9][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N12
cycloneive_lcell_comb \Mux22~13 (
// Equation(s):
// \Mux22~13_combout  = (temp_imemload_output_21 & ((\Mux22~12_combout  & (\storeregister[11][9]~q )) # (!\Mux22~12_combout  & ((\storeregister[9][9]~q ))))) # (!temp_imemload_output_21 & (\Mux22~12_combout ))

	.dataa(temp_imemload_output_21),
	.datab(\Mux22~12_combout ),
	.datac(\storeregister[11][9]~q ),
	.datad(\storeregister[9][9]~q ),
	.cin(gnd),
	.combout(\Mux22~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~13 .lut_mask = 16'hE6C4;
defparam \Mux22~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N7
dffeas \storeregister[2][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][9] .is_wysiwyg = "true";
defparam \storeregister[2][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N17
dffeas \storeregister[3][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][9] .is_wysiwyg = "true";
defparam \storeregister[3][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N16
cycloneive_lcell_comb \Mux22~14 (
// Equation(s):
// \Mux22~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][9]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][9]~q ))))

	.dataa(\storeregister[1][9]~q ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[3][9]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux22~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~14 .lut_mask = 16'hC088;
defparam \Mux22~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N6
cycloneive_lcell_comb \Mux22~15 (
// Equation(s):
// \Mux22~15_combout  = (\Mux22~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][9]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][9]~q ),
	.datad(\Mux22~14_combout ),
	.cin(gnd),
	.combout(\Mux22~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~15 .lut_mask = 16'hFF40;
defparam \Mux22~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N24
cycloneive_lcell_comb \Mux22~16 (
// Equation(s):
// \Mux22~16_combout  = (temp_imemload_output_24 & ((\Mux22~13_combout ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((!temp_imemload_output_23 & \Mux22~15_combout ))))

	.dataa(\Mux22~13_combout ),
	.datab(temp_imemload_output_24),
	.datac(temp_imemload_output_23),
	.datad(\Mux22~15_combout ),
	.cin(gnd),
	.combout(\Mux22~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~16 .lut_mask = 16'hCBC8;
defparam \Mux22~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N16
cycloneive_lcell_comb \Mux59~7 (
// Equation(s):
// \Mux59~7_combout  = (temp_imemload_output_19 & ((\storeregister[27][4]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\storeregister[19][4]~q  & !temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[27][4]~q ),
	.datac(\storeregister[19][4]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux59~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~7 .lut_mask = 16'hAAD8;
defparam \Mux59~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N24
cycloneive_lcell_comb \Mux59~8 (
// Equation(s):
// \Mux59~8_combout  = (\Mux59~7_combout  & ((\storeregister[31][4]~q ) # ((!temp_imemload_output_18)))) # (!\Mux59~7_combout  & (((\storeregister[23][4]~q  & temp_imemload_output_18))))

	.dataa(\Mux59~7_combout ),
	.datab(\storeregister[31][4]~q ),
	.datac(\storeregister[23][4]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux59~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~8 .lut_mask = 16'hD8AA;
defparam \Mux59~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N6
cycloneive_lcell_comb \Mux59~0 (
// Equation(s):
// \Mux59~0_combout  = (temp_imemload_output_19 & (((\storeregister[25][4]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[17][4]~q  & ((!temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[17][4]~q ),
	.datac(\storeregister[25][4]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~0 .lut_mask = 16'hAAE4;
defparam \Mux59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N26
cycloneive_lcell_comb \Mux59~1 (
// Equation(s):
// \Mux59~1_combout  = (temp_imemload_output_18 & ((\Mux59~0_combout  & (\storeregister[29][4]~q )) # (!\Mux59~0_combout  & ((\storeregister[21][4]~q ))))) # (!temp_imemload_output_18 & (((\Mux59~0_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[29][4]~q ),
	.datac(\storeregister[21][4]~q ),
	.datad(\Mux59~0_combout ),
	.cin(gnd),
	.combout(\Mux59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~1 .lut_mask = 16'hDDA0;
defparam \Mux59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N0
cycloneive_lcell_comb \Mux59~5 (
// Equation(s):
// \Mux59~5_combout  = (\Mux59~4_combout  & (((\storeregister[28][4]~q )) # (!temp_imemload_output_19))) # (!\Mux59~4_combout  & (temp_imemload_output_19 & ((\storeregister[24][4]~q ))))

	.dataa(\Mux59~4_combout ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[28][4]~q ),
	.datad(\storeregister[24][4]~q ),
	.cin(gnd),
	.combout(\Mux59~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~5 .lut_mask = 16'hE6A2;
defparam \Mux59~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N16
cycloneive_lcell_comb \Mux59~3 (
// Equation(s):
// \Mux59~3_combout  = (\Mux59~2_combout  & ((\storeregister[30][4]~q ) # ((!temp_imemload_output_19)))) # (!\Mux59~2_combout  & (((\storeregister[26][4]~q  & temp_imemload_output_19))))

	.dataa(\Mux59~2_combout ),
	.datab(\storeregister[30][4]~q ),
	.datac(\storeregister[26][4]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux59~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~3 .lut_mask = 16'hD8AA;
defparam \Mux59~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N24
cycloneive_lcell_comb \Mux59~6 (
// Equation(s):
// \Mux59~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\Mux59~3_combout ))) # (!temp_imemload_output_17 & (\Mux59~5_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux59~5_combout ),
	.datac(temp_imemload_output_17),
	.datad(\Mux59~3_combout ),
	.cin(gnd),
	.combout(\Mux59~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~6 .lut_mask = 16'hF4A4;
defparam \Mux59~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N22
cycloneive_lcell_comb \Mux59~13 (
// Equation(s):
// \Mux59~13_combout  = (\Mux59~12_combout  & (((\storeregister[11][4]~q ) # (!temp_imemload_output_16)))) # (!\Mux59~12_combout  & (\storeregister[9][4]~q  & ((temp_imemload_output_16))))

	.dataa(\Mux59~12_combout ),
	.datab(\storeregister[9][4]~q ),
	.datac(\storeregister[11][4]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux59~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~13 .lut_mask = 16'hE4AA;
defparam \Mux59~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N20
cycloneive_lcell_comb \Mux59~14 (
// Equation(s):
// \Mux59~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[3][4]~q ))) # (!temp_imemload_output_17 & (\storeregister[1][4]~q ))))

	.dataa(\storeregister[1][4]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[3][4]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux59~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~14 .lut_mask = 16'hE200;
defparam \Mux59~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N19
dffeas \storeregister[2][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][4] .is_wysiwyg = "true";
defparam \storeregister[2][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N18
cycloneive_lcell_comb \Mux59~15 (
// Equation(s):
// \Mux59~15_combout  = (\Mux59~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][4]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux59~14_combout ),
	.datac(\storeregister[2][4]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux59~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~15 .lut_mask = 16'hCCEC;
defparam \Mux59~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N26
cycloneive_lcell_comb \Mux59~16 (
// Equation(s):
// \Mux59~16_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\Mux59~13_combout )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & ((\Mux59~15_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\Mux59~13_combout ),
	.datad(\Mux59~15_combout ),
	.cin(gnd),
	.combout(\Mux59~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~16 .lut_mask = 16'hB9A8;
defparam \Mux59~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N22
cycloneive_lcell_comb \Mux59~17 (
// Equation(s):
// \Mux59~17_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[13][4]~q )) # (!temp_imemload_output_16 & ((\storeregister[12][4]~q )))))

	.dataa(\storeregister[13][4]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[12][4]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux59~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~17 .lut_mask = 16'hEE30;
defparam \Mux59~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N18
cycloneive_lcell_comb \Mux59~18 (
// Equation(s):
// \Mux59~18_combout  = (temp_imemload_output_17 & ((\Mux59~17_combout  & ((\storeregister[15][4]~q ))) # (!\Mux59~17_combout  & (\storeregister[14][4]~q )))) # (!temp_imemload_output_17 & (((\Mux59~17_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[14][4]~q ),
	.datac(\Mux59~17_combout ),
	.datad(\storeregister[15][4]~q ),
	.cin(gnd),
	.combout(\Mux59~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~18 .lut_mask = 16'hF858;
defparam \Mux59~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N12
cycloneive_lcell_comb \Mux59~10 (
// Equation(s):
// \Mux59~10_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[5][4]~q ))) # (!temp_imemload_output_16 & (\storeregister[4][4]~q ))))

	.dataa(\storeregister[4][4]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][4]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux59~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~10 .lut_mask = 16'hFC22;
defparam \Mux59~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N4
cycloneive_lcell_comb \storeregister[6][4]~feeder (
// Equation(s):
// \storeregister[6][4]~feeder_combout  = Mux27

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux27),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[6][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[6][4]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[6][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y42_N5
dffeas \storeregister[6][4] (
	.clk(!CLK),
	.d(\storeregister[6][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][4] .is_wysiwyg = "true";
defparam \storeregister[6][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N30
cycloneive_lcell_comb \Mux59~11 (
// Equation(s):
// \Mux59~11_combout  = (\Mux59~10_combout  & (((\storeregister[7][4]~q )) # (!temp_imemload_output_17))) # (!\Mux59~10_combout  & (temp_imemload_output_17 & (\storeregister[6][4]~q )))

	.dataa(\Mux59~10_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[6][4]~q ),
	.datad(\storeregister[7][4]~q ),
	.cin(gnd),
	.combout(\Mux59~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~11 .lut_mask = 16'hEA62;
defparam \Mux59~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N24
cycloneive_lcell_comb \storeregister[27][31]~feeder (
// Equation(s):
// \storeregister[27][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux0),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][31]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y36_N25
dffeas \storeregister[27][31] (
	.clk(!CLK),
	.d(\storeregister[27][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][31] .is_wysiwyg = "true";
defparam \storeregister[27][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N21
dffeas \storeregister[19][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][31] .is_wysiwyg = "true";
defparam \storeregister[19][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N20
cycloneive_lcell_comb \Mux0~7 (
// Equation(s):
// \Mux0~7_combout  = (temp_imemload_output_24 & ((\storeregister[27][31]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[19][31]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[27][31]~q ),
	.datac(\storeregister[19][31]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~7 .lut_mask = 16'hAAD8;
defparam \Mux0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N11
dffeas \storeregister[31][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][31] .is_wysiwyg = "true";
defparam \storeregister[31][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N12
cycloneive_lcell_comb \storeregister[23][31]~feeder (
// Equation(s):
// \storeregister[23][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux0),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[23][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][31]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[23][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N13
dffeas \storeregister[23][31] (
	.clk(!CLK),
	.d(\storeregister[23][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][31] .is_wysiwyg = "true";
defparam \storeregister[23][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N10
cycloneive_lcell_comb \Mux0~8 (
// Equation(s):
// \Mux0~8_combout  = (\Mux0~7_combout  & (((\storeregister[31][31]~q )) # (!temp_imemload_output_23))) # (!\Mux0~7_combout  & (temp_imemload_output_23 & ((\storeregister[23][31]~q ))))

	.dataa(\Mux0~7_combout ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[31][31]~q ),
	.datad(\storeregister[23][31]~q ),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~8 .lut_mask = 16'hE6A2;
defparam \Mux0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N28
cycloneive_lcell_comb \storeregister[26][31]~feeder (
// Equation(s):
// \storeregister[26][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux0),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[26][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[26][31]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[26][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N29
dffeas \storeregister[26][31] (
	.clk(!CLK),
	.d(\storeregister[26][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][31] .is_wysiwyg = "true";
defparam \storeregister[26][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N12
cycloneive_lcell_comb \storeregister[30][31]~feeder (
// Equation(s):
// \storeregister[30][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux0),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[30][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][31]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[30][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N13
dffeas \storeregister[30][31] (
	.clk(!CLK),
	.d(\storeregister[30][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][31] .is_wysiwyg = "true";
defparam \storeregister[30][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N10
cycloneive_lcell_comb \Mux0~3 (
// Equation(s):
// \Mux0~3_combout  = (\Mux0~2_combout  & (((\storeregister[30][31]~q ) # (!temp_imemload_output_24)))) # (!\Mux0~2_combout  & (\storeregister[26][31]~q  & (temp_imemload_output_24)))

	.dataa(\Mux0~2_combout ),
	.datab(\storeregister[26][31]~q ),
	.datac(temp_imemload_output_24),
	.datad(\storeregister[30][31]~q ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~3 .lut_mask = 16'hEA4A;
defparam \Mux0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N3
dffeas \storeregister[20][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][31] .is_wysiwyg = "true";
defparam \storeregister[20][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N2
cycloneive_lcell_comb \Mux0~4 (
// Equation(s):
// \Mux0~4_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[20][31]~q ))) # (!temp_imemload_output_23 & (\storeregister[16][31]~q ))))

	.dataa(\storeregister[16][31]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[20][31]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~4 .lut_mask = 16'hFC22;
defparam \Mux0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N28
cycloneive_lcell_comb \storeregister[24][31]~feeder (
// Equation(s):
// \storeregister[24][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux0),
	.cin(gnd),
	.combout(\storeregister[24][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][31]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[24][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N29
dffeas \storeregister[24][31] (
	.clk(!CLK),
	.d(\storeregister[24][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][31] .is_wysiwyg = "true";
defparam \storeregister[24][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N20
cycloneive_lcell_comb \Mux0~5 (
// Equation(s):
// \Mux0~5_combout  = (temp_imemload_output_24 & ((\Mux0~4_combout  & (\storeregister[28][31]~q )) # (!\Mux0~4_combout  & ((\storeregister[24][31]~q ))))) # (!temp_imemload_output_24 & (((\Mux0~4_combout ))))

	.dataa(\storeregister[28][31]~q ),
	.datab(temp_imemload_output_24),
	.datac(\Mux0~4_combout ),
	.datad(\storeregister[24][31]~q ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~5 .lut_mask = 16'hBCB0;
defparam \Mux0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N24
cycloneive_lcell_comb \Mux0~6 (
// Equation(s):
// \Mux0~6_combout  = (temp_imemload_output_22 & ((\Mux0~3_combout ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((\Mux0~5_combout  & !temp_imemload_output_21))))

	.dataa(\Mux0~3_combout ),
	.datab(\Mux0~5_combout ),
	.datac(temp_imemload_output_22),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~6 .lut_mask = 16'hF0AC;
defparam \Mux0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N3
dffeas \storeregister[25][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][31] .is_wysiwyg = "true";
defparam \storeregister[25][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N2
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (temp_imemload_output_24 & (((\storeregister[25][31]~q ) # (temp_imemload_output_23)))) # (!temp_imemload_output_24 & (\storeregister[17][31]~q  & ((!temp_imemload_output_23))))

	.dataa(\storeregister[17][31]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[25][31]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hCCE2;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N13
dffeas \storeregister[21][31] (
	.clk(!CLK),
	.d(Mux0),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][31] .is_wysiwyg = "true";
defparam \storeregister[21][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N3
dffeas \storeregister[29][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][31] .is_wysiwyg = "true";
defparam \storeregister[29][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N2
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (\Mux0~0_combout  & (((\storeregister[29][31]~q ) # (!temp_imemload_output_23)))) # (!\Mux0~0_combout  & (\storeregister[21][31]~q  & ((temp_imemload_output_23))))

	.dataa(\Mux0~0_combout ),
	.datab(\storeregister[21][31]~q ),
	.datac(\storeregister[29][31]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hE4AA;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N22
cycloneive_lcell_comb \storeregister[15][31]~feeder (
// Equation(s):
// \storeregister[15][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux0),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[15][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][31]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[15][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N23
dffeas \storeregister[15][31] (
	.clk(!CLK),
	.d(\storeregister[15][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][31] .is_wysiwyg = "true";
defparam \storeregister[15][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N31
dffeas \storeregister[14][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][31] .is_wysiwyg = "true";
defparam \storeregister[14][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N25
dffeas \storeregister[12][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][31] .is_wysiwyg = "true";
defparam \storeregister[12][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N28
cycloneive_lcell_comb \Mux0~17 (
// Equation(s):
// \Mux0~17_combout  = (temp_imemload_output_21 & ((\storeregister[13][31]~q ) # ((temp_imemload_output_22)))) # (!temp_imemload_output_21 & (((\storeregister[12][31]~q  & !temp_imemload_output_22))))

	.dataa(\storeregister[13][31]~q ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[12][31]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~17 .lut_mask = 16'hCCB8;
defparam \Mux0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N30
cycloneive_lcell_comb \Mux0~18 (
// Equation(s):
// \Mux0~18_combout  = (temp_imemload_output_22 & ((\Mux0~17_combout  & (\storeregister[15][31]~q )) # (!\Mux0~17_combout  & ((\storeregister[14][31]~q ))))) # (!temp_imemload_output_22 & (((\Mux0~17_combout ))))

	.dataa(\storeregister[15][31]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[14][31]~q ),
	.datad(\Mux0~17_combout ),
	.cin(gnd),
	.combout(\Mux0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~18 .lut_mask = 16'hBBC0;
defparam \Mux0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N29
dffeas \storeregister[2][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][31] .is_wysiwyg = "true";
defparam \storeregister[2][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N5
dffeas \storeregister[3][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][31] .is_wysiwyg = "true";
defparam \storeregister[3][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N4
cycloneive_lcell_comb \Mux0~14 (
// Equation(s):
// \Mux0~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][31]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][31]~q ))))

	.dataa(\storeregister[1][31]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[3][31]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~14 .lut_mask = 16'hE200;
defparam \Mux0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N28
cycloneive_lcell_comb \Mux0~15 (
// Equation(s):
// \Mux0~15_combout  = (\Mux0~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][31]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][31]~q ),
	.datad(\Mux0~14_combout ),
	.cin(gnd),
	.combout(\Mux0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~15 .lut_mask = 16'hFF40;
defparam \Mux0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N20
cycloneive_lcell_comb \storeregister[9][31]~feeder (
// Equation(s):
// \storeregister[9][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux0),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[9][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[9][31]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[9][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N21
dffeas \storeregister[9][31] (
	.clk(!CLK),
	.d(\storeregister[9][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][31] .is_wysiwyg = "true";
defparam \storeregister[9][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N7
dffeas \storeregister[11][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][31] .is_wysiwyg = "true";
defparam \storeregister[11][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N6
cycloneive_lcell_comb \Mux0~13 (
// Equation(s):
// \Mux0~13_combout  = (\Mux0~12_combout  & (((\storeregister[11][31]~q ) # (!temp_imemload_output_21)))) # (!\Mux0~12_combout  & (\storeregister[9][31]~q  & ((temp_imemload_output_21))))

	.dataa(\Mux0~12_combout ),
	.datab(\storeregister[9][31]~q ),
	.datac(\storeregister[11][31]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~13 .lut_mask = 16'hE4AA;
defparam \Mux0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N0
cycloneive_lcell_comb \Mux0~16 (
// Equation(s):
// \Mux0~16_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\Mux0~13_combout ))) # (!temp_imemload_output_24 & (\Mux0~15_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\Mux0~15_combout ),
	.datad(\Mux0~13_combout ),
	.cin(gnd),
	.combout(\Mux0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~16 .lut_mask = 16'hDC98;
defparam \Mux0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y40_N5
dffeas \storeregister[5][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][31] .is_wysiwyg = "true";
defparam \storeregister[5][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N19
dffeas \storeregister[4][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][31] .is_wysiwyg = "true";
defparam \storeregister[4][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N4
cycloneive_lcell_comb \Mux0~10 (
// Equation(s):
// \Mux0~10_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[5][31]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[4][31]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[5][31]~q ),
	.datad(\storeregister[4][31]~q ),
	.cin(gnd),
	.combout(\Mux0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~10 .lut_mask = 16'hB9A8;
defparam \Mux0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N11
dffeas \storeregister[6][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][31] .is_wysiwyg = "true";
defparam \storeregister[6][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N17
dffeas \storeregister[7][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][31] .is_wysiwyg = "true";
defparam \storeregister[7][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N10
cycloneive_lcell_comb \Mux0~11 (
// Equation(s):
// \Mux0~11_combout  = (\Mux0~10_combout  & (((\storeregister[7][31]~q )) # (!temp_imemload_output_22))) # (!\Mux0~10_combout  & (temp_imemload_output_22 & (\storeregister[6][31]~q )))

	.dataa(\Mux0~10_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[6][31]~q ),
	.datad(\storeregister[7][31]~q ),
	.cin(gnd),
	.combout(\Mux0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~11 .lut_mask = 16'hEA62;
defparam \Mux0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N3
dffeas \storeregister[29][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][30] .is_wysiwyg = "true";
defparam \storeregister[29][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N15
dffeas \storeregister[21][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][30] .is_wysiwyg = "true";
defparam \storeregister[21][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N4
cycloneive_lcell_comb \storeregister[17][30]~feeder (
// Equation(s):
// \storeregister[17][30]~feeder_combout  = Mux1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux1),
	.cin(gnd),
	.combout(\storeregister[17][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[17][30]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[17][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N5
dffeas \storeregister[17][30] (
	.clk(!CLK),
	.d(\storeregister[17][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][30] .is_wysiwyg = "true";
defparam \storeregister[17][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N14
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[21][30]~q )) # (!temp_imemload_output_23 & ((\storeregister[17][30]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[21][30]~q ),
	.datad(\storeregister[17][30]~q ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hD9C8;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N13
dffeas \storeregister[25][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][30] .is_wysiwyg = "true";
defparam \storeregister[25][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N2
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (temp_imemload_output_24 & ((\Mux1~0_combout  & (\storeregister[29][30]~q )) # (!\Mux1~0_combout  & ((\storeregister[25][30]~q ))))) # (!temp_imemload_output_24 & (((\Mux1~0_combout ))))

	.dataa(\storeregister[29][30]~q ),
	.datab(temp_imemload_output_24),
	.datac(\Mux1~0_combout ),
	.datad(\storeregister[25][30]~q ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hBCB0;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N19
dffeas \storeregister[30][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][30] .is_wysiwyg = "true";
defparam \storeregister[30][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N29
dffeas \storeregister[26][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][30] .is_wysiwyg = "true";
defparam \storeregister[26][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N28
cycloneive_lcell_comb \Mux1~2 (
// Equation(s):
// \Mux1~2_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[26][30]~q ))) # (!temp_imemload_output_24 & (\storeregister[18][30]~q ))))

	.dataa(\storeregister[18][30]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[26][30]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~2 .lut_mask = 16'hFC22;
defparam \Mux1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N14
cycloneive_lcell_comb \Mux1~3 (
// Equation(s):
// \Mux1~3_combout  = (temp_imemload_output_23 & ((\Mux1~2_combout  & ((\storeregister[30][30]~q ))) # (!\Mux1~2_combout  & (\storeregister[22][30]~q )))) # (!temp_imemload_output_23 & (((\Mux1~2_combout ))))

	.dataa(\storeregister[22][30]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[30][30]~q ),
	.datad(\Mux1~2_combout ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~3 .lut_mask = 16'hF388;
defparam \Mux1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N3
dffeas \storeregister[20][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][30] .is_wysiwyg = "true";
defparam \storeregister[20][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N29
dffeas \storeregister[28][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][30] .is_wysiwyg = "true";
defparam \storeregister[28][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y35_N9
dffeas \storeregister[16][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][30] .is_wysiwyg = "true";
defparam \storeregister[16][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N11
dffeas \storeregister[24][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][30] .is_wysiwyg = "true";
defparam \storeregister[24][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N8
cycloneive_lcell_comb \Mux1~4 (
// Equation(s):
// \Mux1~4_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[24][30]~q ))) # (!temp_imemload_output_24 & (\storeregister[16][30]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][30]~q ),
	.datad(\storeregister[24][30]~q ),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~4 .lut_mask = 16'hDC98;
defparam \Mux1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N28
cycloneive_lcell_comb \Mux1~5 (
// Equation(s):
// \Mux1~5_combout  = (temp_imemload_output_23 & ((\Mux1~4_combout  & ((\storeregister[28][30]~q ))) # (!\Mux1~4_combout  & (\storeregister[20][30]~q )))) # (!temp_imemload_output_23 & (((\Mux1~4_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[20][30]~q ),
	.datac(\storeregister[28][30]~q ),
	.datad(\Mux1~4_combout ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~5 .lut_mask = 16'hF588;
defparam \Mux1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N20
cycloneive_lcell_comb \Mux1~6 (
// Equation(s):
// \Mux1~6_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22)))) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\Mux1~3_combout )) # (!temp_imemload_output_22 & ((\Mux1~5_combout )))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux1~3_combout ),
	.datac(temp_imemload_output_22),
	.datad(\Mux1~5_combout ),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~6 .lut_mask = 16'hE5E0;
defparam \Mux1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N25
dffeas \storeregister[23][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][30] .is_wysiwyg = "true";
defparam \storeregister[23][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N1
dffeas \storeregister[19][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][30] .is_wysiwyg = "true";
defparam \storeregister[19][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N0
cycloneive_lcell_comb \Mux1~7 (
// Equation(s):
// \Mux1~7_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[23][30]~q )) # (!temp_imemload_output_23 & ((\storeregister[19][30]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[23][30]~q ),
	.datac(\storeregister[19][30]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~7 .lut_mask = 16'hEE50;
defparam \Mux1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N31
dffeas \storeregister[31][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][30] .is_wysiwyg = "true";
defparam \storeregister[31][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N27
dffeas \storeregister[27][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][30] .is_wysiwyg = "true";
defparam \storeregister[27][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N30
cycloneive_lcell_comb \Mux1~8 (
// Equation(s):
// \Mux1~8_combout  = (\Mux1~7_combout  & (((\storeregister[31][30]~q )) # (!temp_imemload_output_24))) # (!\Mux1~7_combout  & (temp_imemload_output_24 & ((\storeregister[27][30]~q ))))

	.dataa(\Mux1~7_combout ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[31][30]~q ),
	.datad(\storeregister[27][30]~q ),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~8 .lut_mask = 16'hE6A2;
defparam \Mux1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N26
cycloneive_lcell_comb \storeregister[15][30]~feeder (
// Equation(s):
// \storeregister[15][30]~feeder_combout  = Mux1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux1),
	.cin(gnd),
	.combout(\storeregister[15][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][30]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N27
dffeas \storeregister[15][30] (
	.clk(!CLK),
	.d(\storeregister[15][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][30] .is_wysiwyg = "true";
defparam \storeregister[15][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N24
cycloneive_lcell_comb \storeregister[14][30]~feeder (
// Equation(s):
// \storeregister[14][30]~feeder_combout  = Mux1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux1),
	.cin(gnd),
	.combout(\storeregister[14][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][30]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N25
dffeas \storeregister[14][30] (
	.clk(!CLK),
	.d(\storeregister[14][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][30] .is_wysiwyg = "true";
defparam \storeregister[14][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N11
dffeas \storeregister[13][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][30] .is_wysiwyg = "true";
defparam \storeregister[13][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N15
dffeas \storeregister[12][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][30] .is_wysiwyg = "true";
defparam \storeregister[12][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N14
cycloneive_lcell_comb \Mux1~17 (
// Equation(s):
// \Mux1~17_combout  = (temp_imemload_output_21 & ((\storeregister[13][30]~q ) # ((temp_imemload_output_22)))) # (!temp_imemload_output_21 & (((\storeregister[12][30]~q  & !temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[13][30]~q ),
	.datac(\storeregister[12][30]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux1~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~17 .lut_mask = 16'hAAD8;
defparam \Mux1~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N0
cycloneive_lcell_comb \Mux1~18 (
// Equation(s):
// \Mux1~18_combout  = (\Mux1~17_combout  & ((\storeregister[15][30]~q ) # ((!temp_imemload_output_22)))) # (!\Mux1~17_combout  & (((\storeregister[14][30]~q  & temp_imemload_output_22))))

	.dataa(\storeregister[15][30]~q ),
	.datab(\storeregister[14][30]~q ),
	.datac(\Mux1~17_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux1~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~18 .lut_mask = 16'hACF0;
defparam \Mux1~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N5
dffeas \storeregister[7][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][30] .is_wysiwyg = "true";
defparam \storeregister[7][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y39_N3
dffeas \storeregister[6][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][30] .is_wysiwyg = "true";
defparam \storeregister[6][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N4
cycloneive_lcell_comb \Mux1~13 (
// Equation(s):
// \Mux1~13_combout  = (\Mux1~12_combout  & (((\storeregister[7][30]~q )) # (!temp_imemload_output_22))) # (!\Mux1~12_combout  & (temp_imemload_output_22 & ((\storeregister[6][30]~q ))))

	.dataa(\Mux1~12_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[7][30]~q ),
	.datad(\storeregister[6][30]~q ),
	.cin(gnd),
	.combout(\Mux1~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~13 .lut_mask = 16'hE6A2;
defparam \Mux1~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N17
dffeas \storeregister[2][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][30] .is_wysiwyg = "true";
defparam \storeregister[2][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N15
dffeas \storeregister[1][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][30] .is_wysiwyg = "true";
defparam \storeregister[1][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N25
dffeas \storeregister[3][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][30] .is_wysiwyg = "true";
defparam \storeregister[3][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N24
cycloneive_lcell_comb \Mux1~14 (
// Equation(s):
// \Mux1~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][30]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][30]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[1][30]~q ),
	.datac(\storeregister[3][30]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux1~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~14 .lut_mask = 16'hA088;
defparam \Mux1~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N16
cycloneive_lcell_comb \Mux1~15 (
// Equation(s):
// \Mux1~15_combout  = (\Mux1~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][30]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][30]~q ),
	.datad(\Mux1~14_combout ),
	.cin(gnd),
	.combout(\Mux1~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~15 .lut_mask = 16'hFF40;
defparam \Mux1~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N22
cycloneive_lcell_comb \Mux1~16 (
// Equation(s):
// \Mux1~16_combout  = (temp_imemload_output_23 & ((\Mux1~13_combout ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\Mux1~15_combout  & !temp_imemload_output_24))))

	.dataa(\Mux1~13_combout ),
	.datab(temp_imemload_output_23),
	.datac(\Mux1~15_combout ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux1~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~16 .lut_mask = 16'hCCB8;
defparam \Mux1~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N1
dffeas \storeregister[10][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][30] .is_wysiwyg = "true";
defparam \storeregister[10][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N0
cycloneive_lcell_comb \Mux1~10 (
// Equation(s):
// \Mux1~10_combout  = (temp_imemload_output_22 & (((\storeregister[10][30]~q ) # (temp_imemload_output_21)))) # (!temp_imemload_output_22 & (\storeregister[8][30]~q  & ((!temp_imemload_output_21))))

	.dataa(\storeregister[8][30]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][30]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~10 .lut_mask = 16'hCCE2;
defparam \Mux1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N29
dffeas \storeregister[11][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][30] .is_wysiwyg = "true";
defparam \storeregister[11][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N31
dffeas \storeregister[9][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][30] .is_wysiwyg = "true";
defparam \storeregister[9][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N30
cycloneive_lcell_comb \Mux1~11 (
// Equation(s):
// \Mux1~11_combout  = (\Mux1~10_combout  & ((\storeregister[11][30]~q ) # ((!temp_imemload_output_21)))) # (!\Mux1~10_combout  & (((\storeregister[9][30]~q  & temp_imemload_output_21))))

	.dataa(\Mux1~10_combout ),
	.datab(\storeregister[11][30]~q ),
	.datac(\storeregister[9][30]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux1~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~11 .lut_mask = 16'hD8AA;
defparam \Mux1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N19
dffeas \storeregister[30][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][29] .is_wysiwyg = "true";
defparam \storeregister[30][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N9
dffeas \storeregister[26][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][29] .is_wysiwyg = "true";
defparam \storeregister[26][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N29
dffeas \storeregister[22][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][29] .is_wysiwyg = "true";
defparam \storeregister[22][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N23
dffeas \storeregister[18][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][29] .is_wysiwyg = "true";
defparam \storeregister[18][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N28
cycloneive_lcell_comb \Mux2~2 (
// Equation(s):
// \Mux2~2_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[22][29]~q )) # (!temp_imemload_output_23 & ((\storeregister[18][29]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[22][29]~q ),
	.datad(\storeregister[18][29]~q ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~2 .lut_mask = 16'hD9C8;
defparam \Mux2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N8
cycloneive_lcell_comb \Mux2~3 (
// Equation(s):
// \Mux2~3_combout  = (temp_imemload_output_24 & ((\Mux2~2_combout  & (\storeregister[30][29]~q )) # (!\Mux2~2_combout  & ((\storeregister[26][29]~q ))))) # (!temp_imemload_output_24 & (((\Mux2~2_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[30][29]~q ),
	.datac(\storeregister[26][29]~q ),
	.datad(\Mux2~2_combout ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~3 .lut_mask = 16'hDDA0;
defparam \Mux2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N13
dffeas \storeregister[24][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][29] .is_wysiwyg = "true";
defparam \storeregister[24][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N19
dffeas \storeregister[16][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][29] .is_wysiwyg = "true";
defparam \storeregister[16][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N18
cycloneive_lcell_comb \Mux2~4 (
// Equation(s):
// \Mux2~4_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[20][29]~q )) # (!temp_imemload_output_23 & ((\storeregister[16][29]~q )))))

	.dataa(\storeregister[20][29]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][29]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~4 .lut_mask = 16'hEE30;
defparam \Mux2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N12
cycloneive_lcell_comb \Mux2~5 (
// Equation(s):
// \Mux2~5_combout  = (temp_imemload_output_24 & ((\Mux2~4_combout  & (\storeregister[28][29]~q )) # (!\Mux2~4_combout  & ((\storeregister[24][29]~q ))))) # (!temp_imemload_output_24 & (((\Mux2~4_combout ))))

	.dataa(\storeregister[28][29]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[24][29]~q ),
	.datad(\Mux2~4_combout ),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~5 .lut_mask = 16'hBBC0;
defparam \Mux2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N4
cycloneive_lcell_comb \Mux2~6 (
// Equation(s):
// \Mux2~6_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22)))) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\Mux2~3_combout )) # (!temp_imemload_output_22 & ((\Mux2~5_combout )))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux2~3_combout ),
	.datac(temp_imemload_output_22),
	.datad(\Mux2~5_combout ),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~6 .lut_mask = 16'hE5E0;
defparam \Mux2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N6
cycloneive_lcell_comb \storeregister[29][29]~feeder (
// Equation(s):
// \storeregister[29][29]~feeder_combout  = Mux2

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux2),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[29][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][29]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[29][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N7
dffeas \storeregister[29][29] (
	.clk(!CLK),
	.d(\storeregister[29][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][29] .is_wysiwyg = "true";
defparam \storeregister[29][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N25
dffeas \storeregister[25][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][29] .is_wysiwyg = "true";
defparam \storeregister[25][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N11
dffeas \storeregister[17][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][29] .is_wysiwyg = "true";
defparam \storeregister[17][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N24
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[25][29]~q )) # (!temp_imemload_output_24 & ((\storeregister[17][29]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[25][29]~q ),
	.datad(\storeregister[17][29]~q ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hD9C8;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N0
cycloneive_lcell_comb \storeregister[21][29]~feeder (
// Equation(s):
// \storeregister[21][29]~feeder_combout  = Mux2

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux2),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[21][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][29]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[21][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N1
dffeas \storeregister[21][29] (
	.clk(!CLK),
	.d(\storeregister[21][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][29] .is_wysiwyg = "true";
defparam \storeregister[21][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N18
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (\Mux2~0_combout  & ((\storeregister[29][29]~q ) # ((!temp_imemload_output_23)))) # (!\Mux2~0_combout  & (((temp_imemload_output_23 & \storeregister[21][29]~q ))))

	.dataa(\storeregister[29][29]~q ),
	.datab(\Mux2~0_combout ),
	.datac(temp_imemload_output_23),
	.datad(\storeregister[21][29]~q ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hBC8C;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N15
dffeas \storeregister[27][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][29] .is_wysiwyg = "true";
defparam \storeregister[27][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N19
dffeas \storeregister[19][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][29] .is_wysiwyg = "true";
defparam \storeregister[19][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N18
cycloneive_lcell_comb \Mux2~7 (
// Equation(s):
// \Mux2~7_combout  = (temp_imemload_output_24 & ((\storeregister[27][29]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[19][29]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[27][29]~q ),
	.datac(\storeregister[19][29]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~7 .lut_mask = 16'hAAD8;
defparam \Mux2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N17
dffeas \storeregister[31][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][29] .is_wysiwyg = "true";
defparam \storeregister[31][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N6
cycloneive_lcell_comb \storeregister[23][29]~feeder (
// Equation(s):
// \storeregister[23][29]~feeder_combout  = Mux2

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux2),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[23][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][29]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[23][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N7
dffeas \storeregister[23][29] (
	.clk(!CLK),
	.d(\storeregister[23][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][29] .is_wysiwyg = "true";
defparam \storeregister[23][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N16
cycloneive_lcell_comb \Mux2~8 (
// Equation(s):
// \Mux2~8_combout  = (temp_imemload_output_23 & ((\Mux2~7_combout  & (\storeregister[31][29]~q )) # (!\Mux2~7_combout  & ((\storeregister[23][29]~q ))))) # (!temp_imemload_output_23 & (\Mux2~7_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux2~7_combout ),
	.datac(\storeregister[31][29]~q ),
	.datad(\storeregister[23][29]~q ),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~8 .lut_mask = 16'hE6C4;
defparam \Mux2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N4
cycloneive_lcell_comb \storeregister[12][29]~feeder (
// Equation(s):
// \storeregister[12][29]~feeder_combout  = Mux2

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux2),
	.cin(gnd),
	.combout(\storeregister[12][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[12][29]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[12][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N5
dffeas \storeregister[12][29] (
	.clk(!CLK),
	.d(\storeregister[12][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][29] .is_wysiwyg = "true";
defparam \storeregister[12][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N29
dffeas \storeregister[13][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][29] .is_wysiwyg = "true";
defparam \storeregister[13][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N6
cycloneive_lcell_comb \Mux2~17 (
// Equation(s):
// \Mux2~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][29]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[12][29]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[12][29]~q ),
	.datad(\storeregister[13][29]~q ),
	.cin(gnd),
	.combout(\Mux2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~17 .lut_mask = 16'hBA98;
defparam \Mux2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N31
dffeas \storeregister[14][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][29] .is_wysiwyg = "true";
defparam \storeregister[14][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N28
cycloneive_lcell_comb \storeregister[15][29]~feeder (
// Equation(s):
// \storeregister[15][29]~feeder_combout  = Mux2

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux2),
	.cin(gnd),
	.combout(\storeregister[15][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][29]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y42_N29
dffeas \storeregister[15][29] (
	.clk(!CLK),
	.d(\storeregister[15][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][29] .is_wysiwyg = "true";
defparam \storeregister[15][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N10
cycloneive_lcell_comb \Mux2~18 (
// Equation(s):
// \Mux2~18_combout  = (\Mux2~17_combout  & (((\storeregister[15][29]~q )) # (!temp_imemload_output_22))) # (!\Mux2~17_combout  & (temp_imemload_output_22 & (\storeregister[14][29]~q )))

	.dataa(\Mux2~17_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[14][29]~q ),
	.datad(\storeregister[15][29]~q ),
	.cin(gnd),
	.combout(\Mux2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~18 .lut_mask = 16'hEA62;
defparam \Mux2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N4
cycloneive_lcell_comb \storeregister[9][29]~feeder (
// Equation(s):
// \storeregister[9][29]~feeder_combout  = Mux2

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux2),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[9][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[9][29]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[9][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N5
dffeas \storeregister[9][29] (
	.clk(!CLK),
	.d(\storeregister[9][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][29] .is_wysiwyg = "true";
defparam \storeregister[9][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N11
dffeas \storeregister[11][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][29] .is_wysiwyg = "true";
defparam \storeregister[11][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N9
dffeas \storeregister[10][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][29] .is_wysiwyg = "true";
defparam \storeregister[10][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N23
dffeas \storeregister[8][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][29] .is_wysiwyg = "true";
defparam \storeregister[8][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N22
cycloneive_lcell_comb \Mux2~12 (
// Equation(s):
// \Mux2~12_combout  = (temp_imemload_output_22 & ((\storeregister[10][29]~q ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((\storeregister[8][29]~q  & !temp_imemload_output_21))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[10][29]~q ),
	.datac(\storeregister[8][29]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~12 .lut_mask = 16'hAAD8;
defparam \Mux2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N10
cycloneive_lcell_comb \Mux2~13 (
// Equation(s):
// \Mux2~13_combout  = (temp_imemload_output_21 & ((\Mux2~12_combout  & ((\storeregister[11][29]~q ))) # (!\Mux2~12_combout  & (\storeregister[9][29]~q )))) # (!temp_imemload_output_21 & (((\Mux2~12_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[9][29]~q ),
	.datac(\storeregister[11][29]~q ),
	.datad(\Mux2~12_combout ),
	.cin(gnd),
	.combout(\Mux2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~13 .lut_mask = 16'hF588;
defparam \Mux2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N21
dffeas \storeregister[2][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][29] .is_wysiwyg = "true";
defparam \storeregister[2][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N20
cycloneive_lcell_comb \Mux2~15 (
// Equation(s):
// \Mux2~15_combout  = (\Mux2~14_combout ) # ((temp_imemload_output_22 & (\storeregister[2][29]~q  & !temp_imemload_output_21)))

	.dataa(\Mux2~14_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][29]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~15 .lut_mask = 16'hAAEA;
defparam \Mux2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N30
cycloneive_lcell_comb \Mux2~16 (
// Equation(s):
// \Mux2~16_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\Mux2~13_combout )) # (!temp_imemload_output_24 & ((\Mux2~15_combout )))))

	.dataa(\Mux2~13_combout ),
	.datab(temp_imemload_output_23),
	.datac(temp_imemload_output_24),
	.datad(\Mux2~15_combout ),
	.cin(gnd),
	.combout(\Mux2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~16 .lut_mask = 16'hE3E0;
defparam \Mux2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N23
dffeas \storeregister[7][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][29] .is_wysiwyg = "true";
defparam \storeregister[7][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N13
dffeas \storeregister[6][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][29] .is_wysiwyg = "true";
defparam \storeregister[6][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N21
dffeas \storeregister[5][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][29] .is_wysiwyg = "true";
defparam \storeregister[5][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N3
dffeas \storeregister[4][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][29] .is_wysiwyg = "true";
defparam \storeregister[4][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N20
cycloneive_lcell_comb \Mux2~10 (
// Equation(s):
// \Mux2~10_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[5][29]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[4][29]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[5][29]~q ),
	.datad(\storeregister[4][29]~q ),
	.cin(gnd),
	.combout(\Mux2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~10 .lut_mask = 16'hB9A8;
defparam \Mux2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N12
cycloneive_lcell_comb \Mux2~11 (
// Equation(s):
// \Mux2~11_combout  = (temp_imemload_output_22 & ((\Mux2~10_combout  & (\storeregister[7][29]~q )) # (!\Mux2~10_combout  & ((\storeregister[6][29]~q ))))) # (!temp_imemload_output_22 & (((\Mux2~10_combout ))))

	.dataa(\storeregister[7][29]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[6][29]~q ),
	.datad(\Mux2~10_combout ),
	.cin(gnd),
	.combout(\Mux2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~11 .lut_mask = 16'hBBC0;
defparam \Mux2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N20
cycloneive_lcell_comb \storeregister[23][26]~feeder (
// Equation(s):
// \storeregister[23][26]~feeder_combout  = Mux5

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux5),
	.cin(gnd),
	.combout(\storeregister[23][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][26]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[23][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N21
dffeas \storeregister[23][26] (
	.clk(!CLK),
	.d(\storeregister[23][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][26] .is_wysiwyg = "true";
defparam \storeregister[23][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N9
dffeas \storeregister[19][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][26] .is_wysiwyg = "true";
defparam \storeregister[19][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N8
cycloneive_lcell_comb \Mux5~7 (
// Equation(s):
// \Mux5~7_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[23][26]~q )) # (!temp_imemload_output_23 & ((\storeregister[19][26]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[23][26]~q ),
	.datac(\storeregister[19][26]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~7 .lut_mask = 16'hEE50;
defparam \Mux5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N23
dffeas \storeregister[31][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][26] .is_wysiwyg = "true";
defparam \storeregister[31][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N25
dffeas \storeregister[27][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][26] .is_wysiwyg = "true";
defparam \storeregister[27][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N22
cycloneive_lcell_comb \Mux5~8 (
// Equation(s):
// \Mux5~8_combout  = (temp_imemload_output_24 & ((\Mux5~7_combout  & (\storeregister[31][26]~q )) # (!\Mux5~7_combout  & ((\storeregister[27][26]~q ))))) # (!temp_imemload_output_24 & (\Mux5~7_combout ))

	.dataa(temp_imemload_output_24),
	.datab(\Mux5~7_combout ),
	.datac(\storeregister[31][26]~q ),
	.datad(\storeregister[27][26]~q ),
	.cin(gnd),
	.combout(\Mux5~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~8 .lut_mask = 16'hE6C4;
defparam \Mux5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N21
dffeas \storeregister[16][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][26] .is_wysiwyg = "true";
defparam \storeregister[16][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N19
dffeas \storeregister[24][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][26] .is_wysiwyg = "true";
defparam \storeregister[24][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N20
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[24][26]~q ))) # (!temp_imemload_output_24 & (\storeregister[16][26]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][26]~q ),
	.datad(\storeregister[24][26]~q ),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'hDC98;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N28
cycloneive_lcell_comb \storeregister[28][26]~feeder (
// Equation(s):
// \storeregister[28][26]~feeder_combout  = Mux5

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux5),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[28][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][26]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[28][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N29
dffeas \storeregister[28][26] (
	.clk(!CLK),
	.d(\storeregister[28][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][26] .is_wysiwyg = "true";
defparam \storeregister[28][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N26
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (temp_imemload_output_23 & ((\Mux5~4_combout  & ((\storeregister[28][26]~q ))) # (!\Mux5~4_combout  & (\storeregister[20][26]~q )))) # (!temp_imemload_output_23 & (((\Mux5~4_combout ))))

	.dataa(\storeregister[20][26]~q ),
	.datab(temp_imemload_output_23),
	.datac(\Mux5~4_combout ),
	.datad(\storeregister[28][26]~q ),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'hF838;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N13
dffeas \storeregister[26][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][26] .is_wysiwyg = "true";
defparam \storeregister[26][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N12
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[26][26]~q ))) # (!temp_imemload_output_24 & (\storeregister[18][26]~q ))))

	.dataa(\storeregister[18][26]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[26][26]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'hFC22;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N21
dffeas \storeregister[22][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][26] .is_wysiwyg = "true";
defparam \storeregister[22][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N0
cycloneive_lcell_comb \storeregister[30][26]~feeder (
// Equation(s):
// \storeregister[30][26]~feeder_combout  = Mux5

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux5),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[30][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][26]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[30][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N1
dffeas \storeregister[30][26] (
	.clk(!CLK),
	.d(\storeregister[30][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][26] .is_wysiwyg = "true";
defparam \storeregister[30][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N20
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (temp_imemload_output_23 & ((\Mux5~2_combout  & ((\storeregister[30][26]~q ))) # (!\Mux5~2_combout  & (\storeregister[22][26]~q )))) # (!temp_imemload_output_23 & (\Mux5~2_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux5~2_combout ),
	.datac(\storeregister[22][26]~q ),
	.datad(\storeregister[30][26]~q ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'hEC64;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N14
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// \Mux5~6_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22)))) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & ((\Mux5~3_combout ))) # (!temp_imemload_output_22 & (\Mux5~5_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(\Mux5~5_combout ),
	.datac(\Mux5~3_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'hFA44;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N6
cycloneive_lcell_comb \storeregister[29][26]~feeder (
// Equation(s):
// \storeregister[29][26]~feeder_combout  = Mux5

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux5),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[29][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][26]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[29][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N7
dffeas \storeregister[29][26] (
	.clk(!CLK),
	.d(\storeregister[29][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][26] .is_wysiwyg = "true";
defparam \storeregister[29][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N10
cycloneive_lcell_comb \storeregister[21][26]~feeder (
// Equation(s):
// \storeregister[21][26]~feeder_combout  = Mux5

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux5),
	.cin(gnd),
	.combout(\storeregister[21][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][26]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[21][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N11
dffeas \storeregister[21][26] (
	.clk(!CLK),
	.d(\storeregister[21][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][26] .is_wysiwyg = "true";
defparam \storeregister[21][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N24
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[21][26]~q ))) # (!temp_imemload_output_23 & (\storeregister[17][26]~q ))))

	.dataa(\storeregister[17][26]~q ),
	.datab(temp_imemload_output_24),
	.datac(temp_imemload_output_23),
	.datad(\storeregister[21][26]~q ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hF2C2;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N25
dffeas \storeregister[25][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][26] .is_wysiwyg = "true";
defparam \storeregister[25][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N24
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (\Mux5~0_combout  & ((\storeregister[29][26]~q ) # ((!temp_imemload_output_24)))) # (!\Mux5~0_combout  & (((\storeregister[25][26]~q  & temp_imemload_output_24))))

	.dataa(\storeregister[29][26]~q ),
	.datab(\Mux5~0_combout ),
	.datac(\storeregister[25][26]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hB8CC;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N6
cycloneive_lcell_comb \storeregister[9][26]~feeder (
// Equation(s):
// \storeregister[9][26]~feeder_combout  = Mux5

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux5),
	.cin(gnd),
	.combout(\storeregister[9][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[9][26]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[9][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N7
dffeas \storeregister[9][26] (
	.clk(!CLK),
	.d(\storeregister[9][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][26] .is_wysiwyg = "true";
defparam \storeregister[9][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y41_N23
dffeas \storeregister[11][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][26] .is_wysiwyg = "true";
defparam \storeregister[11][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y39_N7
dffeas \storeregister[10][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][26] .is_wysiwyg = "true";
defparam \storeregister[10][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N6
cycloneive_lcell_comb \Mux5~10 (
// Equation(s):
// \Mux5~10_combout  = (temp_imemload_output_22 & (((\storeregister[10][26]~q ) # (temp_imemload_output_21)))) # (!temp_imemload_output_22 & (\storeregister[8][26]~q  & ((!temp_imemload_output_21))))

	.dataa(\storeregister[8][26]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][26]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux5~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~10 .lut_mask = 16'hCCE2;
defparam \Mux5~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N16
cycloneive_lcell_comb \Mux5~11 (
// Equation(s):
// \Mux5~11_combout  = (temp_imemload_output_21 & ((\Mux5~10_combout  & ((\storeregister[11][26]~q ))) # (!\Mux5~10_combout  & (\storeregister[9][26]~q )))) # (!temp_imemload_output_21 & (((\Mux5~10_combout ))))

	.dataa(\storeregister[9][26]~q ),
	.datab(\storeregister[11][26]~q ),
	.datac(temp_imemload_output_21),
	.datad(\Mux5~10_combout ),
	.cin(gnd),
	.combout(\Mux5~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~11 .lut_mask = 16'hCFA0;
defparam \Mux5~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N11
dffeas \storeregister[14][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][26] .is_wysiwyg = "true";
defparam \storeregister[14][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N16
cycloneive_lcell_comb \storeregister[15][26]~feeder (
// Equation(s):
// \storeregister[15][26]~feeder_combout  = Mux5

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux5),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[15][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][26]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[15][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N17
dffeas \storeregister[15][26] (
	.clk(!CLK),
	.d(\storeregister[15][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][26] .is_wysiwyg = "true";
defparam \storeregister[15][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N1
dffeas \storeregister[13][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][26] .is_wysiwyg = "true";
defparam \storeregister[13][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N31
dffeas \storeregister[12][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][26] .is_wysiwyg = "true";
defparam \storeregister[12][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N30
cycloneive_lcell_comb \Mux5~17 (
// Equation(s):
// \Mux5~17_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & (\storeregister[13][26]~q )) # (!temp_imemload_output_21 & ((\storeregister[12][26]~q )))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[13][26]~q ),
	.datac(\storeregister[12][26]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux5~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~17 .lut_mask = 16'hEE50;
defparam \Mux5~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N30
cycloneive_lcell_comb \Mux5~18 (
// Equation(s):
// \Mux5~18_combout  = (\Mux5~17_combout  & (((\storeregister[15][26]~q ) # (!temp_imemload_output_22)))) # (!\Mux5~17_combout  & (\storeregister[14][26]~q  & ((temp_imemload_output_22))))

	.dataa(\storeregister[14][26]~q ),
	.datab(\storeregister[15][26]~q ),
	.datac(\Mux5~17_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux5~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~18 .lut_mask = 16'hCAF0;
defparam \Mux5~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N25
dffeas \storeregister[2][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][26] .is_wysiwyg = "true";
defparam \storeregister[2][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N21
dffeas \storeregister[3][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][26] .is_wysiwyg = "true";
defparam \storeregister[3][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N20
cycloneive_lcell_comb \Mux5~14 (
// Equation(s):
// \Mux5~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][26]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][26]~q ))))

	.dataa(\storeregister[1][26]~q ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[3][26]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux5~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~14 .lut_mask = 16'hC088;
defparam \Mux5~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N24
cycloneive_lcell_comb \Mux5~15 (
// Equation(s):
// \Mux5~15_combout  = (\Mux5~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][26]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][26]~q ),
	.datad(\Mux5~14_combout ),
	.cin(gnd),
	.combout(\Mux5~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~15 .lut_mask = 16'hFF40;
defparam \Mux5~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N27
dffeas \storeregister[7][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][26] .is_wysiwyg = "true";
defparam \storeregister[7][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N1
dffeas \storeregister[6][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][26] .is_wysiwyg = "true";
defparam \storeregister[6][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N26
cycloneive_lcell_comb \Mux5~13 (
// Equation(s):
// \Mux5~13_combout  = (\Mux5~12_combout  & (((\storeregister[7][26]~q )) # (!temp_imemload_output_22))) # (!\Mux5~12_combout  & (temp_imemload_output_22 & ((\storeregister[6][26]~q ))))

	.dataa(\Mux5~12_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[7][26]~q ),
	.datad(\storeregister[6][26]~q ),
	.cin(gnd),
	.combout(\Mux5~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~13 .lut_mask = 16'hE6A2;
defparam \Mux5~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N24
cycloneive_lcell_comb \Mux5~16 (
// Equation(s):
// \Mux5~16_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\Mux5~13_combout ))) # (!temp_imemload_output_23 & (\Mux5~15_combout ))))

	.dataa(\Mux5~15_combout ),
	.datab(\Mux5~13_combout ),
	.datac(temp_imemload_output_24),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux5~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~16 .lut_mask = 16'hFC0A;
defparam \Mux5~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N24
cycloneive_lcell_comb \storeregister[30][25]~feeder (
// Equation(s):
// \storeregister[30][25]~feeder_combout  = Mux6

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux6),
	.cin(gnd),
	.combout(\storeregister[30][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][25]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[30][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N25
dffeas \storeregister[30][25] (
	.clk(!CLK),
	.d(\storeregister[30][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][25] .is_wysiwyg = "true";
defparam \storeregister[30][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N15
dffeas \storeregister[18][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][25] .is_wysiwyg = "true";
defparam \storeregister[18][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N27
dffeas \storeregister[22][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][25] .is_wysiwyg = "true";
defparam \storeregister[22][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N26
cycloneive_lcell_comb \Mux6~2 (
// Equation(s):
// \Mux6~2_combout  = (temp_imemload_output_23 & (((\storeregister[22][25]~q ) # (temp_imemload_output_24)))) # (!temp_imemload_output_23 & (\storeregister[18][25]~q  & ((!temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[18][25]~q ),
	.datac(\storeregister[22][25]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~2 .lut_mask = 16'hAAE4;
defparam \Mux6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N14
cycloneive_lcell_comb \Mux6~3 (
// Equation(s):
// \Mux6~3_combout  = (temp_imemload_output_24 & ((\Mux6~2_combout  & ((\storeregister[30][25]~q ))) # (!\Mux6~2_combout  & (\storeregister[26][25]~q )))) # (!temp_imemload_output_24 & (((\Mux6~2_combout ))))

	.dataa(\storeregister[26][25]~q ),
	.datab(\storeregister[30][25]~q ),
	.datac(temp_imemload_output_24),
	.datad(\Mux6~2_combout ),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~3 .lut_mask = 16'hCFA0;
defparam \Mux6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N15
dffeas \storeregister[16][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][25] .is_wysiwyg = "true";
defparam \storeregister[16][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N12
cycloneive_lcell_comb \storeregister[20][25]~feeder (
// Equation(s):
// \storeregister[20][25]~feeder_combout  = Mux6

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux6),
	.cin(gnd),
	.combout(\storeregister[20][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][25]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[20][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N13
dffeas \storeregister[20][25] (
	.clk(!CLK),
	.d(\storeregister[20][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][25] .is_wysiwyg = "true";
defparam \storeregister[20][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N14
cycloneive_lcell_comb \Mux6~4 (
// Equation(s):
// \Mux6~4_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[20][25]~q ))) # (!temp_imemload_output_23 & (\storeregister[16][25]~q ))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[16][25]~q ),
	.datad(\storeregister[20][25]~q ),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~4 .lut_mask = 16'hDC98;
defparam \Mux6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N23
dffeas \storeregister[28][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][25] .is_wysiwyg = "true";
defparam \storeregister[28][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N22
cycloneive_lcell_comb \Mux6~5 (
// Equation(s):
// \Mux6~5_combout  = (\Mux6~4_combout  & (((\storeregister[28][25]~q ) # (!temp_imemload_output_24)))) # (!\Mux6~4_combout  & (\storeregister[24][25]~q  & ((temp_imemload_output_24))))

	.dataa(\storeregister[24][25]~q ),
	.datab(\Mux6~4_combout ),
	.datac(\storeregister[28][25]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~5 .lut_mask = 16'hE2CC;
defparam \Mux6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N30
cycloneive_lcell_comb \Mux6~6 (
// Equation(s):
// \Mux6~6_combout  = (temp_imemload_output_22 & ((\Mux6~3_combout ) # ((temp_imemload_output_21)))) # (!temp_imemload_output_22 & (((!temp_imemload_output_21 & \Mux6~5_combout ))))

	.dataa(\Mux6~3_combout ),
	.datab(temp_imemload_output_22),
	.datac(temp_imemload_output_21),
	.datad(\Mux6~5_combout ),
	.cin(gnd),
	.combout(\Mux6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~6 .lut_mask = 16'hCBC8;
defparam \Mux6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N9
dffeas \storeregister[31][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][25] .is_wysiwyg = "true";
defparam \storeregister[31][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N30
cycloneive_lcell_comb \storeregister[19][25]~feeder (
// Equation(s):
// \storeregister[19][25]~feeder_combout  = Mux6

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux6),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[19][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[19][25]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[19][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N31
dffeas \storeregister[19][25] (
	.clk(!CLK),
	.d(\storeregister[19][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][25] .is_wysiwyg = "true";
defparam \storeregister[19][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N21
dffeas \storeregister[27][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][25] .is_wysiwyg = "true";
defparam \storeregister[27][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N20
cycloneive_lcell_comb \Mux6~7 (
// Equation(s):
// \Mux6~7_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[27][25]~q ))) # (!temp_imemload_output_24 & (\storeregister[19][25]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[19][25]~q ),
	.datac(\storeregister[27][25]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux6~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~7 .lut_mask = 16'hFA44;
defparam \Mux6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N11
dffeas \storeregister[23][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][25] .is_wysiwyg = "true";
defparam \storeregister[23][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N8
cycloneive_lcell_comb \Mux6~8 (
// Equation(s):
// \Mux6~8_combout  = (\Mux6~7_combout  & ((\storeregister[31][25]~q ) # ((!temp_imemload_output_23)))) # (!\Mux6~7_combout  & (((\storeregister[23][25]~q  & temp_imemload_output_23))))

	.dataa(\storeregister[31][25]~q ),
	.datab(\Mux6~7_combout ),
	.datac(\storeregister[23][25]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux6~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~8 .lut_mask = 16'hB8CC;
defparam \Mux6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N8
cycloneive_lcell_comb \storeregister[29][25]~feeder (
// Equation(s):
// \storeregister[29][25]~feeder_combout  = Mux6

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux6),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[29][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[29][25]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[29][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N9
dffeas \storeregister[29][25] (
	.clk(!CLK),
	.d(\storeregister[29][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][25] .is_wysiwyg = "true";
defparam \storeregister[29][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N0
cycloneive_lcell_comb \storeregister[21][25]~feeder (
// Equation(s):
// \storeregister[21][25]~feeder_combout  = Mux6

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux6),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[21][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][25]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[21][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N1
dffeas \storeregister[21][25] (
	.clk(!CLK),
	.d(\storeregister[21][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][25] .is_wysiwyg = "true";
defparam \storeregister[21][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N15
dffeas \storeregister[25][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][25] .is_wysiwyg = "true";
defparam \storeregister[25][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N22
cycloneive_lcell_comb \storeregister[17][25]~feeder (
// Equation(s):
// \storeregister[17][25]~feeder_combout  = Mux6

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux6),
	.cin(gnd),
	.combout(\storeregister[17][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[17][25]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[17][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N23
dffeas \storeregister[17][25] (
	.clk(!CLK),
	.d(\storeregister[17][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][25] .is_wysiwyg = "true";
defparam \storeregister[17][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N14
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[25][25]~q )) # (!temp_imemload_output_24 & ((\storeregister[17][25]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[25][25]~q ),
	.datad(\storeregister[17][25]~q ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hD9C8;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N28
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (\Mux6~0_combout  & ((\storeregister[29][25]~q ) # ((!temp_imemload_output_23)))) # (!\Mux6~0_combout  & (((\storeregister[21][25]~q  & temp_imemload_output_23))))

	.dataa(\storeregister[29][25]~q ),
	.datab(\storeregister[21][25]~q ),
	.datac(\Mux6~0_combout ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hACF0;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N4
cycloneive_lcell_comb \storeregister[15][25]~feeder (
// Equation(s):
// \storeregister[15][25]~feeder_combout  = Mux6

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux6),
	.cin(gnd),
	.combout(\storeregister[15][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][25]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N5
dffeas \storeregister[15][25] (
	.clk(!CLK),
	.d(\storeregister[15][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][25] .is_wysiwyg = "true";
defparam \storeregister[15][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N3
dffeas \storeregister[12][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][25] .is_wysiwyg = "true";
defparam \storeregister[12][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N25
dffeas \storeregister[13][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][25] .is_wysiwyg = "true";
defparam \storeregister[13][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N2
cycloneive_lcell_comb \Mux6~17 (
// Equation(s):
// \Mux6~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][25]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[12][25]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[12][25]~q ),
	.datad(\storeregister[13][25]~q ),
	.cin(gnd),
	.combout(\Mux6~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~17 .lut_mask = 16'hBA98;
defparam \Mux6~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N1
dffeas \storeregister[14][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][25] .is_wysiwyg = "true";
defparam \storeregister[14][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N22
cycloneive_lcell_comb \Mux6~18 (
// Equation(s):
// \Mux6~18_combout  = (temp_imemload_output_22 & ((\Mux6~17_combout  & (\storeregister[15][25]~q )) # (!\Mux6~17_combout  & ((\storeregister[14][25]~q ))))) # (!temp_imemload_output_22 & (((\Mux6~17_combout ))))

	.dataa(\storeregister[15][25]~q ),
	.datab(temp_imemload_output_22),
	.datac(\Mux6~17_combout ),
	.datad(\storeregister[14][25]~q ),
	.cin(gnd),
	.combout(\Mux6~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~18 .lut_mask = 16'hBCB0;
defparam \Mux6~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N29
dffeas \storeregister[9][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][25] .is_wysiwyg = "true";
defparam \storeregister[9][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N3
dffeas \storeregister[11][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][25] .is_wysiwyg = "true";
defparam \storeregister[11][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N2
cycloneive_lcell_comb \Mux6~13 (
// Equation(s):
// \Mux6~13_combout  = (\Mux6~12_combout  & (((\storeregister[11][25]~q ) # (!temp_imemload_output_21)))) # (!\Mux6~12_combout  & (\storeregister[9][25]~q  & ((temp_imemload_output_21))))

	.dataa(\Mux6~12_combout ),
	.datab(\storeregister[9][25]~q ),
	.datac(\storeregister[11][25]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux6~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~13 .lut_mask = 16'hE4AA;
defparam \Mux6~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N1
dffeas \storeregister[2][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][25] .is_wysiwyg = "true";
defparam \storeregister[2][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N9
dffeas \storeregister[3][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][25] .is_wysiwyg = "true";
defparam \storeregister[3][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N8
cycloneive_lcell_comb \Mux6~14 (
// Equation(s):
// \Mux6~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][25]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][25]~q ))))

	.dataa(\storeregister[1][25]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[3][25]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux6~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~14 .lut_mask = 16'hE200;
defparam \Mux6~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N0
cycloneive_lcell_comb \Mux6~15 (
// Equation(s):
// \Mux6~15_combout  = (\Mux6~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][25]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][25]~q ),
	.datad(\Mux6~14_combout ),
	.cin(gnd),
	.combout(\Mux6~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~15 .lut_mask = 16'hFF40;
defparam \Mux6~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N8
cycloneive_lcell_comb \Mux6~16 (
// Equation(s):
// \Mux6~16_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\Mux6~13_combout )) # (!temp_imemload_output_24 & ((\Mux6~15_combout )))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\Mux6~13_combout ),
	.datad(\Mux6~15_combout ),
	.cin(gnd),
	.combout(\Mux6~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~16 .lut_mask = 16'hD9C8;
defparam \Mux6~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N7
dffeas \storeregister[7][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][25] .is_wysiwyg = "true";
defparam \storeregister[7][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N21
dffeas \storeregister[6][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][25] .is_wysiwyg = "true";
defparam \storeregister[6][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y41_N5
dffeas \storeregister[5][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][25] .is_wysiwyg = "true";
defparam \storeregister[5][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N4
cycloneive_lcell_comb \Mux6~10 (
// Equation(s):
// \Mux6~10_combout  = (temp_imemload_output_21 & (((\storeregister[5][25]~q ) # (temp_imemload_output_22)))) # (!temp_imemload_output_21 & (\storeregister[4][25]~q  & ((!temp_imemload_output_22))))

	.dataa(\storeregister[4][25]~q ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[5][25]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux6~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~10 .lut_mask = 16'hCCE2;
defparam \Mux6~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N20
cycloneive_lcell_comb \Mux6~11 (
// Equation(s):
// \Mux6~11_combout  = (temp_imemload_output_22 & ((\Mux6~10_combout  & (\storeregister[7][25]~q )) # (!\Mux6~10_combout  & ((\storeregister[6][25]~q ))))) # (!temp_imemload_output_22 & (((\Mux6~10_combout ))))

	.dataa(\storeregister[7][25]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[6][25]~q ),
	.datad(\Mux6~10_combout ),
	.cin(gnd),
	.combout(\Mux6~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~11 .lut_mask = 16'hBBC0;
defparam \Mux6~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N11
dffeas \storeregister[20][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][28] .is_wysiwyg = "true";
defparam \storeregister[20][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N0
cycloneive_lcell_comb \storeregister[16][28]~feeder (
// Equation(s):
// \storeregister[16][28]~feeder_combout  = Mux3

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux3),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[16][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[16][28]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[16][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N1
dffeas \storeregister[16][28] (
	.clk(!CLK),
	.d(\storeregister[16][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][28] .is_wysiwyg = "true";
defparam \storeregister[16][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N0
cycloneive_lcell_comb \storeregister[24][28]~feeder (
// Equation(s):
// \storeregister[24][28]~feeder_combout  = Mux3

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux3),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[24][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][28]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[24][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N1
dffeas \storeregister[24][28] (
	.clk(!CLK),
	.d(\storeregister[24][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][28] .is_wysiwyg = "true";
defparam \storeregister[24][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N2
cycloneive_lcell_comb \Mux3~4 (
// Equation(s):
// \Mux3~4_combout  = (temp_imemload_output_24 & ((temp_imemload_output_23) # ((\storeregister[24][28]~q )))) # (!temp_imemload_output_24 & (!temp_imemload_output_23 & (\storeregister[16][28]~q )))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[16][28]~q ),
	.datad(\storeregister[24][28]~q ),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~4 .lut_mask = 16'hBA98;
defparam \Mux3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N6
cycloneive_lcell_comb \Mux3~5 (
// Equation(s):
// \Mux3~5_combout  = (temp_imemload_output_23 & ((\Mux3~4_combout  & (\storeregister[28][28]~q )) # (!\Mux3~4_combout  & ((\storeregister[20][28]~q ))))) # (!temp_imemload_output_23 & (((\Mux3~4_combout ))))

	.dataa(\storeregister[28][28]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[20][28]~q ),
	.datad(\Mux3~4_combout ),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~5 .lut_mask = 16'hBBC0;
defparam \Mux3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N26
cycloneive_lcell_comb \storeregister[30][28]~feeder (
// Equation(s):
// \storeregister[30][28]~feeder_combout  = Mux3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux3),
	.cin(gnd),
	.combout(\storeregister[30][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][28]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[30][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N27
dffeas \storeregister[30][28] (
	.clk(!CLK),
	.d(\storeregister[30][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][28] .is_wysiwyg = "true";
defparam \storeregister[30][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N21
dffeas \storeregister[26][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][28] .is_wysiwyg = "true";
defparam \storeregister[26][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N20
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[26][28]~q ))) # (!temp_imemload_output_24 & (\storeregister[18][28]~q ))))

	.dataa(\storeregister[18][28]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[26][28]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hFC22;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N12
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// \Mux3~3_combout  = (temp_imemload_output_23 & ((\Mux3~2_combout  & ((\storeregister[30][28]~q ))) # (!\Mux3~2_combout  & (\storeregister[22][28]~q )))) # (!temp_imemload_output_23 & (((\Mux3~2_combout ))))

	.dataa(\storeregister[22][28]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[30][28]~q ),
	.datad(\Mux3~2_combout ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hF388;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N20
cycloneive_lcell_comb \Mux3~6 (
// Equation(s):
// \Mux3~6_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22)))) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & ((\Mux3~3_combout ))) # (!temp_imemload_output_22 & (\Mux3~5_combout ))))

	.dataa(\Mux3~5_combout ),
	.datab(\Mux3~3_combout ),
	.datac(temp_imemload_output_21),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~6 .lut_mask = 16'hFC0A;
defparam \Mux3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N9
dffeas \storeregister[31][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][28] .is_wysiwyg = "true";
defparam \storeregister[31][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N14
cycloneive_lcell_comb \storeregister[19][28]~feeder (
// Equation(s):
// \storeregister[19][28]~feeder_combout  = Mux3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux3),
	.cin(gnd),
	.combout(\storeregister[19][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[19][28]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[19][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N15
dffeas \storeregister[19][28] (
	.clk(!CLK),
	.d(\storeregister[19][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][28] .is_wysiwyg = "true";
defparam \storeregister[19][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N5
dffeas \storeregister[23][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][28] .is_wysiwyg = "true";
defparam \storeregister[23][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N4
cycloneive_lcell_comb \Mux3~7 (
// Equation(s):
// \Mux3~7_combout  = (temp_imemload_output_23 & (((\storeregister[23][28]~q ) # (temp_imemload_output_24)))) # (!temp_imemload_output_23 & (\storeregister[19][28]~q  & ((!temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[19][28]~q ),
	.datac(\storeregister[23][28]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~7 .lut_mask = 16'hAAE4;
defparam \Mux3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N3
dffeas \storeregister[27][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][28] .is_wysiwyg = "true";
defparam \storeregister[27][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N26
cycloneive_lcell_comb \Mux3~8 (
// Equation(s):
// \Mux3~8_combout  = (\Mux3~7_combout  & ((\storeregister[31][28]~q ) # ((!temp_imemload_output_24)))) # (!\Mux3~7_combout  & (((temp_imemload_output_24 & \storeregister[27][28]~q ))))

	.dataa(\storeregister[31][28]~q ),
	.datab(\Mux3~7_combout ),
	.datac(temp_imemload_output_24),
	.datad(\storeregister[27][28]~q ),
	.cin(gnd),
	.combout(\Mux3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~8 .lut_mask = 16'hBC8C;
defparam \Mux3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N9
dffeas \storeregister[25][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][28] .is_wysiwyg = "true";
defparam \storeregister[25][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N15
dffeas \storeregister[29][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][28] .is_wysiwyg = "true";
defparam \storeregister[29][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N28
cycloneive_lcell_comb \storeregister[21][28]~feeder (
// Equation(s):
// \storeregister[21][28]~feeder_combout  = Mux3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux3),
	.cin(gnd),
	.combout(\storeregister[21][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][28]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[21][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N29
dffeas \storeregister[21][28] (
	.clk(!CLK),
	.d(\storeregister[21][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][28] .is_wysiwyg = "true";
defparam \storeregister[21][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N9
dffeas \storeregister[17][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][28] .is_wysiwyg = "true";
defparam \storeregister[17][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N8
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (temp_imemload_output_23 & ((\storeregister[21][28]~q ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\storeregister[17][28]~q  & !temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[21][28]~q ),
	.datac(\storeregister[17][28]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hAAD8;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N14
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (temp_imemload_output_24 & ((\Mux3~0_combout  & ((\storeregister[29][28]~q ))) # (!\Mux3~0_combout  & (\storeregister[25][28]~q )))) # (!temp_imemload_output_24 & (((\Mux3~0_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[25][28]~q ),
	.datac(\storeregister[29][28]~q ),
	.datad(\Mux3~0_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hF588;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N23
dffeas \storeregister[10][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][28] .is_wysiwyg = "true";
defparam \storeregister[10][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N22
cycloneive_lcell_comb \Mux3~10 (
// Equation(s):
// \Mux3~10_combout  = (temp_imemload_output_22 & (((\storeregister[10][28]~q ) # (temp_imemload_output_21)))) # (!temp_imemload_output_22 & (\storeregister[8][28]~q  & ((!temp_imemload_output_21))))

	.dataa(\storeregister[8][28]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][28]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~10 .lut_mask = 16'hCCE2;
defparam \Mux3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N5
dffeas \storeregister[9][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][28] .is_wysiwyg = "true";
defparam \storeregister[9][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N11
dffeas \storeregister[11][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][28] .is_wysiwyg = "true";
defparam \storeregister[11][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N4
cycloneive_lcell_comb \Mux3~11 (
// Equation(s):
// \Mux3~11_combout  = (\Mux3~10_combout  & (((\storeregister[11][28]~q )) # (!temp_imemload_output_21))) # (!\Mux3~10_combout  & (temp_imemload_output_21 & (\storeregister[9][28]~q )))

	.dataa(\Mux3~10_combout ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[9][28]~q ),
	.datad(\storeregister[11][28]~q ),
	.cin(gnd),
	.combout(\Mux3~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~11 .lut_mask = 16'hEA62;
defparam \Mux3~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y40_N15
dffeas \storeregister[15][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][28] .is_wysiwyg = "true";
defparam \storeregister[15][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N24
cycloneive_lcell_comb \storeregister[12][28]~feeder (
// Equation(s):
// \storeregister[12][28]~feeder_combout  = Mux3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux3),
	.cin(gnd),
	.combout(\storeregister[12][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[12][28]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[12][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y40_N25
dffeas \storeregister[12][28] (
	.clk(!CLK),
	.d(\storeregister[12][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][28] .is_wysiwyg = "true";
defparam \storeregister[12][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y40_N12
cycloneive_lcell_comb \storeregister[13][28]~feeder (
// Equation(s):
// \storeregister[13][28]~feeder_combout  = Mux3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux3),
	.cin(gnd),
	.combout(\storeregister[13][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[13][28]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[13][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y40_N13
dffeas \storeregister[13][28] (
	.clk(!CLK),
	.d(\storeregister[13][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][28] .is_wysiwyg = "true";
defparam \storeregister[13][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y40_N2
cycloneive_lcell_comb \Mux3~17 (
// Equation(s):
// \Mux3~17_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22) # (\storeregister[13][28]~q )))) # (!temp_imemload_output_21 & (\storeregister[12][28]~q  & (!temp_imemload_output_22)))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[12][28]~q ),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[13][28]~q ),
	.cin(gnd),
	.combout(\Mux3~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~17 .lut_mask = 16'hAEA4;
defparam \Mux3~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y40_N10
cycloneive_lcell_comb \storeregister[14][28]~feeder (
// Equation(s):
// \storeregister[14][28]~feeder_combout  = Mux3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux3),
	.cin(gnd),
	.combout(\storeregister[14][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][28]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y40_N11
dffeas \storeregister[14][28] (
	.clk(!CLK),
	.d(\storeregister[14][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][28] .is_wysiwyg = "true";
defparam \storeregister[14][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y40_N20
cycloneive_lcell_comb \Mux3~18 (
// Equation(s):
// \Mux3~18_combout  = (\Mux3~17_combout  & ((\storeregister[15][28]~q ) # ((!temp_imemload_output_22)))) # (!\Mux3~17_combout  & (((temp_imemload_output_22 & \storeregister[14][28]~q ))))

	.dataa(\storeregister[15][28]~q ),
	.datab(\Mux3~17_combout ),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[14][28]~q ),
	.cin(gnd),
	.combout(\Mux3~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~18 .lut_mask = 16'hBC8C;
defparam \Mux3~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N31
dffeas \storeregister[2][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][28] .is_wysiwyg = "true";
defparam \storeregister[2][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N13
dffeas \storeregister[3][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][28] .is_wysiwyg = "true";
defparam \storeregister[3][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N12
cycloneive_lcell_comb \Mux3~14 (
// Equation(s):
// \Mux3~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][28]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][28]~q ))))

	.dataa(\storeregister[1][28]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[3][28]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux3~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~14 .lut_mask = 16'hE200;
defparam \Mux3~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N30
cycloneive_lcell_comb \Mux3~15 (
// Equation(s):
// \Mux3~15_combout  = (\Mux3~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][28]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][28]~q ),
	.datad(\Mux3~14_combout ),
	.cin(gnd),
	.combout(\Mux3~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~15 .lut_mask = 16'hFF40;
defparam \Mux3~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N31
dffeas \storeregister[7][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][28] .is_wysiwyg = "true";
defparam \storeregister[7][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N25
dffeas \storeregister[6][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][28] .is_wysiwyg = "true";
defparam \storeregister[6][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N30
cycloneive_lcell_comb \Mux3~13 (
// Equation(s):
// \Mux3~13_combout  = (\Mux3~12_combout  & (((\storeregister[7][28]~q )) # (!temp_imemload_output_22))) # (!\Mux3~12_combout  & (temp_imemload_output_22 & ((\storeregister[6][28]~q ))))

	.dataa(\Mux3~12_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[7][28]~q ),
	.datad(\storeregister[6][28]~q ),
	.cin(gnd),
	.combout(\Mux3~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~13 .lut_mask = 16'hE6A2;
defparam \Mux3~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y40_N0
cycloneive_lcell_comb \Mux3~16 (
// Equation(s):
// \Mux3~16_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\Mux3~13_combout ))) # (!temp_imemload_output_23 & (\Mux3~15_combout ))))

	.dataa(\Mux3~15_combout ),
	.datab(\Mux3~13_combout ),
	.datac(temp_imemload_output_24),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux3~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~16 .lut_mask = 16'hFC0A;
defparam \Mux3~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N1
dffeas \storeregister[27][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][27] .is_wysiwyg = "true";
defparam \storeregister[27][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N9
dffeas \storeregister[19][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][27] .is_wysiwyg = "true";
defparam \storeregister[19][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N8
cycloneive_lcell_comb \Mux4~7 (
// Equation(s):
// \Mux4~7_combout  = (temp_imemload_output_24 & ((\storeregister[27][27]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[19][27]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[27][27]~q ),
	.datac(\storeregister[19][27]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~7 .lut_mask = 16'hAAD8;
defparam \Mux4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N23
dffeas \storeregister[23][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][27] .is_wysiwyg = "true";
defparam \storeregister[23][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N4
cycloneive_lcell_comb \storeregister[31][27]~feeder (
// Equation(s):
// \storeregister[31][27]~feeder_combout  = Mux4

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux4),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[31][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][27]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[31][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N5
dffeas \storeregister[31][27] (
	.clk(!CLK),
	.d(\storeregister[31][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][27] .is_wysiwyg = "true";
defparam \storeregister[31][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N22
cycloneive_lcell_comb \Mux4~8 (
// Equation(s):
// \Mux4~8_combout  = (temp_imemload_output_23 & ((\Mux4~7_combout  & ((\storeregister[31][27]~q ))) # (!\Mux4~7_combout  & (\storeregister[23][27]~q )))) # (!temp_imemload_output_23 & (\Mux4~7_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux4~7_combout ),
	.datac(\storeregister[23][27]~q ),
	.datad(\storeregister[31][27]~q ),
	.cin(gnd),
	.combout(\Mux4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~8 .lut_mask = 16'hEC64;
defparam \Mux4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N29
dffeas \storeregister[25][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][27] .is_wysiwyg = "true";
defparam \storeregister[25][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N11
dffeas \storeregister[17][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][27] .is_wysiwyg = "true";
defparam \storeregister[17][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N10
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (temp_imemload_output_24 & ((\storeregister[25][27]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[17][27]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[25][27]~q ),
	.datac(\storeregister[17][27]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hAAD8;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N19
dffeas \storeregister[29][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][27] .is_wysiwyg = "true";
defparam \storeregister[29][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N2
cycloneive_lcell_comb \storeregister[21][27]~feeder (
// Equation(s):
// \storeregister[21][27]~feeder_combout  = Mux4

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux4),
	.cin(gnd),
	.combout(\storeregister[21][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][27]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[21][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N3
dffeas \storeregister[21][27] (
	.clk(!CLK),
	.d(\storeregister[21][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][27] .is_wysiwyg = "true";
defparam \storeregister[21][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N28
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (\Mux4~0_combout  & ((\storeregister[29][27]~q ) # ((!temp_imemload_output_23)))) # (!\Mux4~0_combout  & (((temp_imemload_output_23 & \storeregister[21][27]~q ))))

	.dataa(\Mux4~0_combout ),
	.datab(\storeregister[29][27]~q ),
	.datac(temp_imemload_output_23),
	.datad(\storeregister[21][27]~q ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hDA8A;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N1
dffeas \storeregister[26][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][27] .is_wysiwyg = "true";
defparam \storeregister[26][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N11
dffeas \storeregister[30][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][27] .is_wysiwyg = "true";
defparam \storeregister[30][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N10
cycloneive_lcell_comb \Mux4~3 (
// Equation(s):
// \Mux4~3_combout  = (\Mux4~2_combout  & (((\storeregister[30][27]~q ) # (!temp_imemload_output_24)))) # (!\Mux4~2_combout  & (\storeregister[26][27]~q  & ((temp_imemload_output_24))))

	.dataa(\Mux4~2_combout ),
	.datab(\storeregister[26][27]~q ),
	.datac(\storeregister[30][27]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~3 .lut_mask = 16'hE4AA;
defparam \Mux4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N21
dffeas \storeregister[20][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][27] .is_wysiwyg = "true";
defparam \storeregister[20][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N7
dffeas \storeregister[16][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][27] .is_wysiwyg = "true";
defparam \storeregister[16][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N20
cycloneive_lcell_comb \Mux4~4 (
// Equation(s):
// \Mux4~4_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\storeregister[20][27]~q )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & ((\storeregister[16][27]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[20][27]~q ),
	.datad(\storeregister[16][27]~q ),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~4 .lut_mask = 16'hB9A8;
defparam \Mux4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N19
dffeas \storeregister[28][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][27] .is_wysiwyg = "true";
defparam \storeregister[28][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N18
cycloneive_lcell_comb \Mux4~5 (
// Equation(s):
// \Mux4~5_combout  = (\Mux4~4_combout  & (((\storeregister[28][27]~q ) # (!temp_imemload_output_24)))) # (!\Mux4~4_combout  & (\storeregister[24][27]~q  & ((temp_imemload_output_24))))

	.dataa(\storeregister[24][27]~q ),
	.datab(\Mux4~4_combout ),
	.datac(\storeregister[28][27]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~5 .lut_mask = 16'hE2CC;
defparam \Mux4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N12
cycloneive_lcell_comb \Mux4~6 (
// Equation(s):
// \Mux4~6_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\Mux4~3_combout )) # (!temp_imemload_output_22 & ((\Mux4~5_combout )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\Mux4~3_combout ),
	.datad(\Mux4~5_combout ),
	.cin(gnd),
	.combout(\Mux4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~6 .lut_mask = 16'hD9C8;
defparam \Mux4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N5
dffeas \storeregister[6][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][27] .is_wysiwyg = "true";
defparam \storeregister[6][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N3
dffeas \storeregister[7][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][27] .is_wysiwyg = "true";
defparam \storeregister[7][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N9
dffeas \storeregister[5][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][27] .is_wysiwyg = "true";
defparam \storeregister[5][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N15
dffeas \storeregister[4][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][27] .is_wysiwyg = "true";
defparam \storeregister[4][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N8
cycloneive_lcell_comb \Mux4~10 (
// Equation(s):
// \Mux4~10_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[5][27]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[4][27]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[5][27]~q ),
	.datad(\storeregister[4][27]~q ),
	.cin(gnd),
	.combout(\Mux4~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~10 .lut_mask = 16'hB9A8;
defparam \Mux4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N2
cycloneive_lcell_comb \Mux4~11 (
// Equation(s):
// \Mux4~11_combout  = (temp_imemload_output_22 & ((\Mux4~10_combout  & ((\storeregister[7][27]~q ))) # (!\Mux4~10_combout  & (\storeregister[6][27]~q )))) # (!temp_imemload_output_22 & (((\Mux4~10_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[6][27]~q ),
	.datac(\storeregister[7][27]~q ),
	.datad(\Mux4~10_combout ),
	.cin(gnd),
	.combout(\Mux4~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~11 .lut_mask = 16'hF588;
defparam \Mux4~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N15
dffeas \storeregister[10][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][27] .is_wysiwyg = "true";
defparam \storeregister[10][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N29
dffeas \storeregister[8][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][27] .is_wysiwyg = "true";
defparam \storeregister[8][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N14
cycloneive_lcell_comb \Mux4~12 (
// Equation(s):
// \Mux4~12_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\storeregister[10][27]~q )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & ((\storeregister[8][27]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[10][27]~q ),
	.datad(\storeregister[8][27]~q ),
	.cin(gnd),
	.combout(\Mux4~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~12 .lut_mask = 16'hB9A8;
defparam \Mux4~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N7
dffeas \storeregister[11][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][27] .is_wysiwyg = "true";
defparam \storeregister[11][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N6
cycloneive_lcell_comb \Mux4~13 (
// Equation(s):
// \Mux4~13_combout  = (\Mux4~12_combout  & (((\storeregister[11][27]~q ) # (!temp_imemload_output_21)))) # (!\Mux4~12_combout  & (\storeregister[9][27]~q  & ((temp_imemload_output_21))))

	.dataa(\storeregister[9][27]~q ),
	.datab(\Mux4~12_combout ),
	.datac(\storeregister[11][27]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux4~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~13 .lut_mask = 16'hE2CC;
defparam \Mux4~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N11
dffeas \storeregister[1][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][27] .is_wysiwyg = "true";
defparam \storeregister[1][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N9
dffeas \storeregister[3][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][27] .is_wysiwyg = "true";
defparam \storeregister[3][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N8
cycloneive_lcell_comb \Mux4~14 (
// Equation(s):
// \Mux4~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][27]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][27]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[1][27]~q ),
	.datac(\storeregister[3][27]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux4~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~14 .lut_mask = 16'hA088;
defparam \Mux4~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N13
dffeas \storeregister[2][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][27] .is_wysiwyg = "true";
defparam \storeregister[2][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N12
cycloneive_lcell_comb \Mux4~15 (
// Equation(s):
// \Mux4~15_combout  = (\Mux4~14_combout ) # ((!temp_imemload_output_21 & (\storeregister[2][27]~q  & temp_imemload_output_22)))

	.dataa(temp_imemload_output_21),
	.datab(\Mux4~14_combout ),
	.datac(\storeregister[2][27]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux4~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~15 .lut_mask = 16'hDCCC;
defparam \Mux4~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N2
cycloneive_lcell_comb \Mux4~16 (
// Equation(s):
// \Mux4~16_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\Mux4~13_combout )) # (!temp_imemload_output_24 & ((\Mux4~15_combout )))))

	.dataa(\Mux4~13_combout ),
	.datab(temp_imemload_output_23),
	.datac(temp_imemload_output_24),
	.datad(\Mux4~15_combout ),
	.cin(gnd),
	.combout(\Mux4~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~16 .lut_mask = 16'hE3E0;
defparam \Mux4~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N30
cycloneive_lcell_comb \storeregister[15][27]~feeder (
// Equation(s):
// \storeregister[15][27]~feeder_combout  = Mux4

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux4),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[15][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][27]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[15][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N31
dffeas \storeregister[15][27] (
	.clk(!CLK),
	.d(\storeregister[15][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][27] .is_wysiwyg = "true";
defparam \storeregister[15][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N20
cycloneive_lcell_comb \storeregister[14][27]~feeder (
// Equation(s):
// \storeregister[14][27]~feeder_combout  = Mux4

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux4),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[14][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][27]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[14][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N21
dffeas \storeregister[14][27] (
	.clk(!CLK),
	.d(\storeregister[14][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][27] .is_wysiwyg = "true";
defparam \storeregister[14][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N3
dffeas \storeregister[12][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][27] .is_wysiwyg = "true";
defparam \storeregister[12][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N2
cycloneive_lcell_comb \Mux4~17 (
// Equation(s):
// \Mux4~17_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & (\storeregister[13][27]~q )) # (!temp_imemload_output_21 & ((\storeregister[12][27]~q )))))

	.dataa(\storeregister[13][27]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[12][27]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux4~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~17 .lut_mask = 16'hEE30;
defparam \Mux4~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N28
cycloneive_lcell_comb \Mux4~18 (
// Equation(s):
// \Mux4~18_combout  = (\Mux4~17_combout  & ((\storeregister[15][27]~q ) # ((!temp_imemload_output_22)))) # (!\Mux4~17_combout  & (((\storeregister[14][27]~q  & temp_imemload_output_22))))

	.dataa(\storeregister[15][27]~q ),
	.datab(\storeregister[14][27]~q ),
	.datac(\Mux4~17_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux4~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~18 .lut_mask = 16'hACF0;
defparam \Mux4~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N22
cycloneive_lcell_comb \storeregister[26][17]~feeder (
// Equation(s):
// \storeregister[26][17]~feeder_combout  = Mux14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux14),
	.cin(gnd),
	.combout(\storeregister[26][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[26][17]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[26][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N23
dffeas \storeregister[26][17] (
	.clk(!CLK),
	.d(\storeregister[26][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][17] .is_wysiwyg = "true";
defparam \storeregister[26][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N2
cycloneive_lcell_comb \storeregister[30][17]~feeder (
// Equation(s):
// \storeregister[30][17]~feeder_combout  = Mux14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux14),
	.cin(gnd),
	.combout(\storeregister[30][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][17]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[30][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N3
dffeas \storeregister[30][17] (
	.clk(!CLK),
	.d(\storeregister[30][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][17] .is_wysiwyg = "true";
defparam \storeregister[30][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N28
cycloneive_lcell_comb \Mux14~3 (
// Equation(s):
// \Mux14~3_combout  = (\Mux14~2_combout  & (((\storeregister[30][17]~q ) # (!temp_imemload_output_24)))) # (!\Mux14~2_combout  & (\storeregister[26][17]~q  & (temp_imemload_output_24)))

	.dataa(\Mux14~2_combout ),
	.datab(\storeregister[26][17]~q ),
	.datac(temp_imemload_output_24),
	.datad(\storeregister[30][17]~q ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~3 .lut_mask = 16'hEA4A;
defparam \Mux14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N27
dffeas \storeregister[16][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][17] .is_wysiwyg = "true";
defparam \storeregister[16][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N26
cycloneive_lcell_comb \Mux14~4 (
// Equation(s):
// \Mux14~4_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[20][17]~q )) # (!temp_imemload_output_23 & ((\storeregister[16][17]~q )))))

	.dataa(\storeregister[20][17]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][17]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~4 .lut_mask = 16'hEE30;
defparam \Mux14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N9
dffeas \storeregister[24][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][17] .is_wysiwyg = "true";
defparam \storeregister[24][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N16
cycloneive_lcell_comb \Mux14~5 (
// Equation(s):
// \Mux14~5_combout  = (\Mux14~4_combout  & ((\storeregister[28][17]~q ) # ((!temp_imemload_output_24)))) # (!\Mux14~4_combout  & (((\storeregister[24][17]~q  & temp_imemload_output_24))))

	.dataa(\storeregister[28][17]~q ),
	.datab(\Mux14~4_combout ),
	.datac(\storeregister[24][17]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~5 .lut_mask = 16'hB8CC;
defparam \Mux14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N10
cycloneive_lcell_comb \Mux14~6 (
// Equation(s):
// \Mux14~6_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\Mux14~3_combout )) # (!temp_imemload_output_22 & ((\Mux14~5_combout )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\Mux14~3_combout ),
	.datad(\Mux14~5_combout ),
	.cin(gnd),
	.combout(\Mux14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~6 .lut_mask = 16'hD9C8;
defparam \Mux14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N11
dffeas \storeregister[23][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][17] .is_wysiwyg = "true";
defparam \storeregister[23][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N13
dffeas \storeregister[31][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][17] .is_wysiwyg = "true";
defparam \storeregister[31][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N6
cycloneive_lcell_comb \storeregister[27][17]~feeder (
// Equation(s):
// \storeregister[27][17]~feeder_combout  = Mux14

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux14),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][17]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N7
dffeas \storeregister[27][17] (
	.clk(!CLK),
	.d(\storeregister[27][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][17] .is_wysiwyg = "true";
defparam \storeregister[27][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N1
dffeas \storeregister[19][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][17] .is_wysiwyg = "true";
defparam \storeregister[19][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N0
cycloneive_lcell_comb \Mux14~7 (
// Equation(s):
// \Mux14~7_combout  = (temp_imemload_output_24 & ((\storeregister[27][17]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[19][17]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[27][17]~q ),
	.datac(\storeregister[19][17]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux14~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~7 .lut_mask = 16'hAAD8;
defparam \Mux14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N4
cycloneive_lcell_comb \Mux14~8 (
// Equation(s):
// \Mux14~8_combout  = (\Mux14~7_combout  & (((\storeregister[31][17]~q ) # (!temp_imemload_output_23)))) # (!\Mux14~7_combout  & (\storeregister[23][17]~q  & ((temp_imemload_output_23))))

	.dataa(\storeregister[23][17]~q ),
	.datab(\storeregister[31][17]~q ),
	.datac(\Mux14~7_combout ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux14~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~8 .lut_mask = 16'hCAF0;
defparam \Mux14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N23
dffeas \storeregister[21][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][17] .is_wysiwyg = "true";
defparam \storeregister[21][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N31
dffeas \storeregister[25][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][17] .is_wysiwyg = "true";
defparam \storeregister[25][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N29
dffeas \storeregister[17][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][17] .is_wysiwyg = "true";
defparam \storeregister[17][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N28
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (temp_imemload_output_24 & ((\storeregister[25][17]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[17][17]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[25][17]~q ),
	.datac(\storeregister[17][17]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hAAD8;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N21
dffeas \storeregister[29][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][17] .is_wysiwyg = "true";
defparam \storeregister[29][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N20
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (\Mux14~0_combout  & (((\storeregister[29][17]~q ) # (!temp_imemload_output_23)))) # (!\Mux14~0_combout  & (\storeregister[21][17]~q  & ((temp_imemload_output_23))))

	.dataa(\storeregister[21][17]~q ),
	.datab(\Mux14~0_combout ),
	.datac(\storeregister[29][17]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hE2CC;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N14
cycloneive_lcell_comb \storeregister[14][17]~feeder (
// Equation(s):
// \storeregister[14][17]~feeder_combout  = Mux14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux14),
	.cin(gnd),
	.combout(\storeregister[14][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][17]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N15
dffeas \storeregister[14][17] (
	.clk(!CLK),
	.d(\storeregister[14][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][17] .is_wysiwyg = "true";
defparam \storeregister[14][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N29
dffeas \storeregister[12][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][17] .is_wysiwyg = "true";
defparam \storeregister[12][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N7
dffeas \storeregister[13][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][17] .is_wysiwyg = "true";
defparam \storeregister[13][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N28
cycloneive_lcell_comb \Mux14~17 (
// Equation(s):
// \Mux14~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][17]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[12][17]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[12][17]~q ),
	.datad(\storeregister[13][17]~q ),
	.cin(gnd),
	.combout(\Mux14~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~17 .lut_mask = 16'hBA98;
defparam \Mux14~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N24
cycloneive_lcell_comb \storeregister[15][17]~feeder (
// Equation(s):
// \storeregister[15][17]~feeder_combout  = Mux14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux14),
	.cin(gnd),
	.combout(\storeregister[15][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][17]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y40_N25
dffeas \storeregister[15][17] (
	.clk(!CLK),
	.d(\storeregister[15][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][17] .is_wysiwyg = "true";
defparam \storeregister[15][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N6
cycloneive_lcell_comb \Mux14~18 (
// Equation(s):
// \Mux14~18_combout  = (temp_imemload_output_22 & ((\Mux14~17_combout  & ((\storeregister[15][17]~q ))) # (!\Mux14~17_combout  & (\storeregister[14][17]~q )))) # (!temp_imemload_output_22 & (((\Mux14~17_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[14][17]~q ),
	.datac(\Mux14~17_combout ),
	.datad(\storeregister[15][17]~q ),
	.cin(gnd),
	.combout(\Mux14~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~18 .lut_mask = 16'hF858;
defparam \Mux14~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N23
dffeas \storeregister[2][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][17] .is_wysiwyg = "true";
defparam \storeregister[2][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N31
dffeas \storeregister[1][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][17] .is_wysiwyg = "true";
defparam \storeregister[1][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N17
dffeas \storeregister[3][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][17] .is_wysiwyg = "true";
defparam \storeregister[3][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N16
cycloneive_lcell_comb \Mux14~14 (
// Equation(s):
// \Mux14~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][17]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][17]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[1][17]~q ),
	.datac(\storeregister[3][17]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux14~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~14 .lut_mask = 16'hE400;
defparam \Mux14~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N22
cycloneive_lcell_comb \Mux14~15 (
// Equation(s):
// \Mux14~15_combout  = (\Mux14~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][17]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][17]~q ),
	.datad(\Mux14~14_combout ),
	.cin(gnd),
	.combout(\Mux14~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~15 .lut_mask = 16'hFF40;
defparam \Mux14~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N7
dffeas \storeregister[8][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][17] .is_wysiwyg = "true";
defparam \storeregister[8][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N29
dffeas \storeregister[10][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][17] .is_wysiwyg = "true";
defparam \storeregister[10][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N6
cycloneive_lcell_comb \Mux14~12 (
// Equation(s):
// \Mux14~12_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\storeregister[10][17]~q )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & (\storeregister[8][17]~q )))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[8][17]~q ),
	.datad(\storeregister[10][17]~q ),
	.cin(gnd),
	.combout(\Mux14~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~12 .lut_mask = 16'hBA98;
defparam \Mux14~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N5
dffeas \storeregister[11][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][17] .is_wysiwyg = "true";
defparam \storeregister[11][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N4
cycloneive_lcell_comb \Mux14~13 (
// Equation(s):
// \Mux14~13_combout  = (\Mux14~12_combout  & (((\storeregister[11][17]~q ) # (!temp_imemload_output_21)))) # (!\Mux14~12_combout  & (\storeregister[9][17]~q  & ((temp_imemload_output_21))))

	.dataa(\storeregister[9][17]~q ),
	.datab(\Mux14~12_combout ),
	.datac(\storeregister[11][17]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux14~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~13 .lut_mask = 16'hE2CC;
defparam \Mux14~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N24
cycloneive_lcell_comb \Mux14~16 (
// Equation(s):
// \Mux14~16_combout  = (temp_imemload_output_24 & (((\Mux14~13_combout ) # (temp_imemload_output_23)))) # (!temp_imemload_output_24 & (\Mux14~15_combout  & ((!temp_imemload_output_23))))

	.dataa(\Mux14~15_combout ),
	.datab(temp_imemload_output_24),
	.datac(\Mux14~13_combout ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux14~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~16 .lut_mask = 16'hCCE2;
defparam \Mux14~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y40_N13
dffeas \storeregister[5][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][17] .is_wysiwyg = "true";
defparam \storeregister[5][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N7
dffeas \storeregister[4][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][17] .is_wysiwyg = "true";
defparam \storeregister[4][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N12
cycloneive_lcell_comb \Mux14~10 (
// Equation(s):
// \Mux14~10_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[5][17]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[4][17]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[5][17]~q ),
	.datad(\storeregister[4][17]~q ),
	.cin(gnd),
	.combout(\Mux14~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~10 .lut_mask = 16'hB9A8;
defparam \Mux14~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N29
dffeas \storeregister[6][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][17] .is_wysiwyg = "true";
defparam \storeregister[6][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N19
dffeas \storeregister[7][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][17] .is_wysiwyg = "true";
defparam \storeregister[7][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N28
cycloneive_lcell_comb \Mux14~11 (
// Equation(s):
// \Mux14~11_combout  = (\Mux14~10_combout  & (((\storeregister[7][17]~q )) # (!temp_imemload_output_22))) # (!\Mux14~10_combout  & (temp_imemload_output_22 & (\storeregister[6][17]~q )))

	.dataa(\Mux14~10_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[6][17]~q ),
	.datad(\storeregister[7][17]~q ),
	.cin(gnd),
	.combout(\Mux14~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~11 .lut_mask = 16'hEA62;
defparam \Mux14~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N11
dffeas \storeregister[31][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][20] .is_wysiwyg = "true";
defparam \storeregister[31][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N21
dffeas \storeregister[27][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][20] .is_wysiwyg = "true";
defparam \storeregister[27][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N11
dffeas \storeregister[19][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][20] .is_wysiwyg = "true";
defparam \storeregister[19][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N10
cycloneive_lcell_comb \Mux11~7 (
// Equation(s):
// \Mux11~7_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[23][20]~q )) # (!temp_imemload_output_23 & ((\storeregister[19][20]~q )))))

	.dataa(\storeregister[23][20]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[19][20]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~7 .lut_mask = 16'hEE30;
defparam \Mux11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N8
cycloneive_lcell_comb \Mux11~8 (
// Equation(s):
// \Mux11~8_combout  = (temp_imemload_output_24 & ((\Mux11~7_combout  & (\storeregister[31][20]~q )) # (!\Mux11~7_combout  & ((\storeregister[27][20]~q ))))) # (!temp_imemload_output_24 & (((\Mux11~7_combout ))))

	.dataa(\storeregister[31][20]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[27][20]~q ),
	.datad(\Mux11~7_combout ),
	.cin(gnd),
	.combout(\Mux11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~8 .lut_mask = 16'hBBC0;
defparam \Mux11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N5
dffeas \storeregister[25][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][20] .is_wysiwyg = "true";
defparam \storeregister[25][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N31
dffeas \storeregister[29][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][20] .is_wysiwyg = "true";
defparam \storeregister[29][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N2
cycloneive_lcell_comb \storeregister[21][20]~feeder (
// Equation(s):
// \storeregister[21][20]~feeder_combout  = Mux11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux11),
	.cin(gnd),
	.combout(\storeregister[21][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][20]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[21][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N3
dffeas \storeregister[21][20] (
	.clk(!CLK),
	.d(\storeregister[21][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][20] .is_wysiwyg = "true";
defparam \storeregister[21][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N19
dffeas \storeregister[17][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][20] .is_wysiwyg = "true";
defparam \storeregister[17][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N18
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[21][20]~q )) # (!temp_imemload_output_23 & ((\storeregister[17][20]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[21][20]~q ),
	.datac(\storeregister[17][20]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hEE50;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N30
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (temp_imemload_output_24 & ((\Mux11~0_combout  & ((\storeregister[29][20]~q ))) # (!\Mux11~0_combout  & (\storeregister[25][20]~q )))) # (!temp_imemload_output_24 & (((\Mux11~0_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[25][20]~q ),
	.datac(\storeregister[29][20]~q ),
	.datad(\Mux11~0_combout ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hF588;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N5
dffeas \storeregister[20][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][20] .is_wysiwyg = "true";
defparam \storeregister[20][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N17
dffeas \storeregister[28][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][20] .is_wysiwyg = "true";
defparam \storeregister[28][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N16
cycloneive_lcell_comb \Mux11~5 (
// Equation(s):
// \Mux11~5_combout  = (\Mux11~4_combout  & (((\storeregister[28][20]~q ) # (!temp_imemload_output_23)))) # (!\Mux11~4_combout  & (\storeregister[20][20]~q  & ((temp_imemload_output_23))))

	.dataa(\Mux11~4_combout ),
	.datab(\storeregister[20][20]~q ),
	.datac(\storeregister[28][20]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~5 .lut_mask = 16'hE4AA;
defparam \Mux11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N21
dffeas \storeregister[30][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][20] .is_wysiwyg = "true";
defparam \storeregister[30][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N11
dffeas \storeregister[22][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][20] .is_wysiwyg = "true";
defparam \storeregister[22][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N24
cycloneive_lcell_comb \storeregister[26][20]~feeder (
// Equation(s):
// \storeregister[26][20]~feeder_combout  = Mux11

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux11),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[26][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[26][20]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[26][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N25
dffeas \storeregister[26][20] (
	.clk(!CLK),
	.d(\storeregister[26][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][20] .is_wysiwyg = "true";
defparam \storeregister[26][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N11
dffeas \storeregister[18][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][20] .is_wysiwyg = "true";
defparam \storeregister[18][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N10
cycloneive_lcell_comb \Mux11~2 (
// Equation(s):
// \Mux11~2_combout  = (temp_imemload_output_24 & ((\storeregister[26][20]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[18][20]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[26][20]~q ),
	.datac(\storeregister[18][20]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~2 .lut_mask = 16'hAAD8;
defparam \Mux11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N2
cycloneive_lcell_comb \Mux11~3 (
// Equation(s):
// \Mux11~3_combout  = (temp_imemload_output_23 & ((\Mux11~2_combout  & (\storeregister[30][20]~q )) # (!\Mux11~2_combout  & ((\storeregister[22][20]~q ))))) # (!temp_imemload_output_23 & (((\Mux11~2_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[30][20]~q ),
	.datac(\storeregister[22][20]~q ),
	.datad(\Mux11~2_combout ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~3 .lut_mask = 16'hDDA0;
defparam \Mux11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N10
cycloneive_lcell_comb \Mux11~6 (
// Equation(s):
// \Mux11~6_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & ((\Mux11~3_combout ))) # (!temp_imemload_output_22 & (\Mux11~5_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\Mux11~5_combout ),
	.datad(\Mux11~3_combout ),
	.cin(gnd),
	.combout(\Mux11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~6 .lut_mask = 16'hDC98;
defparam \Mux11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N22
cycloneive_lcell_comb \storeregister[15][20]~feeder (
// Equation(s):
// \storeregister[15][20]~feeder_combout  = Mux11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux11),
	.cin(gnd),
	.combout(\storeregister[15][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][20]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y40_N23
dffeas \storeregister[15][20] (
	.clk(!CLK),
	.d(\storeregister[15][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][20] .is_wysiwyg = "true";
defparam \storeregister[15][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N31
dffeas \storeregister[12][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][20] .is_wysiwyg = "true";
defparam \storeregister[12][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N21
dffeas \storeregister[13][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][20] .is_wysiwyg = "true";
defparam \storeregister[13][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N30
cycloneive_lcell_comb \Mux11~17 (
// Equation(s):
// \Mux11~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][20]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[12][20]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[12][20]~q ),
	.datad(\storeregister[13][20]~q ),
	.cin(gnd),
	.combout(\Mux11~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~17 .lut_mask = 16'hBA98;
defparam \Mux11~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N0
cycloneive_lcell_comb \storeregister[14][20]~feeder (
// Equation(s):
// \storeregister[14][20]~feeder_combout  = Mux11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux11),
	.cin(gnd),
	.combout(\storeregister[14][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][20]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y40_N1
dffeas \storeregister[14][20] (
	.clk(!CLK),
	.d(\storeregister[14][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][20] .is_wysiwyg = "true";
defparam \storeregister[14][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N16
cycloneive_lcell_comb \Mux11~18 (
// Equation(s):
// \Mux11~18_combout  = (\Mux11~17_combout  & ((\storeregister[15][20]~q ) # ((!temp_imemload_output_22)))) # (!\Mux11~17_combout  & (((temp_imemload_output_22 & \storeregister[14][20]~q ))))

	.dataa(\storeregister[15][20]~q ),
	.datab(\Mux11~17_combout ),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[14][20]~q ),
	.cin(gnd),
	.combout(\Mux11~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~18 .lut_mask = 16'hBC8C;
defparam \Mux11~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N29
dffeas \storeregister[2][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][20] .is_wysiwyg = "true";
defparam \storeregister[2][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N28
cycloneive_lcell_comb \Mux11~15 (
// Equation(s):
// \Mux11~15_combout  = (\Mux11~14_combout ) # ((temp_imemload_output_22 & (\storeregister[2][20]~q  & !temp_imemload_output_21)))

	.dataa(\Mux11~14_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][20]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux11~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~15 .lut_mask = 16'hAAEA;
defparam \Mux11~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N9
dffeas \storeregister[6][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][20] .is_wysiwyg = "true";
defparam \storeregister[6][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N11
dffeas \storeregister[7][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][20] .is_wysiwyg = "true";
defparam \storeregister[7][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y41_N9
dffeas \storeregister[5][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][20] .is_wysiwyg = "true";
defparam \storeregister[5][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y41_N7
dffeas \storeregister[4][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][20] .is_wysiwyg = "true";
defparam \storeregister[4][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N6
cycloneive_lcell_comb \Mux11~12 (
// Equation(s):
// \Mux11~12_combout  = (temp_imemload_output_21 & ((\storeregister[5][20]~q ) # ((temp_imemload_output_22)))) # (!temp_imemload_output_21 & (((\storeregister[4][20]~q  & !temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[5][20]~q ),
	.datac(\storeregister[4][20]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux11~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~12 .lut_mask = 16'hAAD8;
defparam \Mux11~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N10
cycloneive_lcell_comb \Mux11~13 (
// Equation(s):
// \Mux11~13_combout  = (temp_imemload_output_22 & ((\Mux11~12_combout  & ((\storeregister[7][20]~q ))) # (!\Mux11~12_combout  & (\storeregister[6][20]~q )))) # (!temp_imemload_output_22 & (((\Mux11~12_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[6][20]~q ),
	.datac(\storeregister[7][20]~q ),
	.datad(\Mux11~12_combout ),
	.cin(gnd),
	.combout(\Mux11~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~13 .lut_mask = 16'hF588;
defparam \Mux11~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N26
cycloneive_lcell_comb \Mux11~16 (
// Equation(s):
// \Mux11~16_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\Mux11~13_combout ))) # (!temp_imemload_output_23 & (\Mux11~15_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\Mux11~15_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux11~13_combout ),
	.cin(gnd),
	.combout(\Mux11~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~16 .lut_mask = 16'hF4A4;
defparam \Mux11~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N9
dffeas \storeregister[8][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][20] .is_wysiwyg = "true";
defparam \storeregister[8][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N3
dffeas \storeregister[10][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][20] .is_wysiwyg = "true";
defparam \storeregister[10][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N2
cycloneive_lcell_comb \Mux11~10 (
// Equation(s):
// \Mux11~10_combout  = (temp_imemload_output_22 & (((\storeregister[10][20]~q ) # (temp_imemload_output_21)))) # (!temp_imemload_output_22 & (\storeregister[8][20]~q  & ((!temp_imemload_output_21))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[8][20]~q ),
	.datac(\storeregister[10][20]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~10 .lut_mask = 16'hAAE4;
defparam \Mux11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N9
dffeas \storeregister[9][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][20] .is_wysiwyg = "true";
defparam \storeregister[9][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N19
dffeas \storeregister[11][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][20] .is_wysiwyg = "true";
defparam \storeregister[11][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N8
cycloneive_lcell_comb \Mux11~11 (
// Equation(s):
// \Mux11~11_combout  = (\Mux11~10_combout  & (((\storeregister[11][20]~q )) # (!temp_imemload_output_21))) # (!\Mux11~10_combout  & (temp_imemload_output_21 & (\storeregister[9][20]~q )))

	.dataa(\Mux11~10_combout ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[9][20]~q ),
	.datad(\storeregister[11][20]~q ),
	.cin(gnd),
	.combout(\Mux11~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~11 .lut_mask = 16'hEA62;
defparam \Mux11~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N21
dffeas \storeregister[30][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][19] .is_wysiwyg = "true";
defparam \storeregister[30][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N21
dffeas \storeregister[22][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][19] .is_wysiwyg = "true";
defparam \storeregister[22][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N7
dffeas \storeregister[18][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][19] .is_wysiwyg = "true";
defparam \storeregister[18][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N20
cycloneive_lcell_comb \Mux12~2 (
// Equation(s):
// \Mux12~2_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[22][19]~q )) # (!temp_imemload_output_23 & ((\storeregister[18][19]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[22][19]~q ),
	.datad(\storeregister[18][19]~q ),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~2 .lut_mask = 16'hD9C8;
defparam \Mux12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N20
cycloneive_lcell_comb \Mux12~3 (
// Equation(s):
// \Mux12~3_combout  = (temp_imemload_output_24 & ((\Mux12~2_combout  & ((\storeregister[30][19]~q ))) # (!\Mux12~2_combout  & (\storeregister[26][19]~q )))) # (!temp_imemload_output_24 & (((\Mux12~2_combout ))))

	.dataa(\storeregister[26][19]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[30][19]~q ),
	.datad(\Mux12~2_combout ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~3 .lut_mask = 16'hF388;
defparam \Mux12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N9
dffeas \storeregister[28][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][19] .is_wysiwyg = "true";
defparam \storeregister[28][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N11
dffeas \storeregister[16][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][19] .is_wysiwyg = "true";
defparam \storeregister[16][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N3
dffeas \storeregister[20][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][19] .is_wysiwyg = "true";
defparam \storeregister[20][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N2
cycloneive_lcell_comb \Mux12~4 (
// Equation(s):
// \Mux12~4_combout  = (temp_imemload_output_23 & (((\storeregister[20][19]~q ) # (temp_imemload_output_24)))) # (!temp_imemload_output_23 & (\storeregister[16][19]~q  & ((!temp_imemload_output_24))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[16][19]~q ),
	.datac(\storeregister[20][19]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~4 .lut_mask = 16'hAAE4;
defparam \Mux12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N8
cycloneive_lcell_comb \Mux12~5 (
// Equation(s):
// \Mux12~5_combout  = (temp_imemload_output_24 & ((\Mux12~4_combout  & ((\storeregister[28][19]~q ))) # (!\Mux12~4_combout  & (\storeregister[24][19]~q )))) # (!temp_imemload_output_24 & (((\Mux12~4_combout ))))

	.dataa(\storeregister[24][19]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[28][19]~q ),
	.datad(\Mux12~4_combout ),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~5 .lut_mask = 16'hF388;
defparam \Mux12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N18
cycloneive_lcell_comb \Mux12~6 (
// Equation(s):
// \Mux12~6_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\Mux12~3_combout )) # (!temp_imemload_output_22 & ((\Mux12~5_combout )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\Mux12~3_combout ),
	.datad(\Mux12~5_combout ),
	.cin(gnd),
	.combout(\Mux12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~6 .lut_mask = 16'hD9C8;
defparam \Mux12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N13
dffeas \storeregister[25][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][19] .is_wysiwyg = "true";
defparam \storeregister[25][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N31
dffeas \storeregister[17][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][19] .is_wysiwyg = "true";
defparam \storeregister[17][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N12
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[25][19]~q )) # (!temp_imemload_output_24 & ((\storeregister[17][19]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[25][19]~q ),
	.datad(\storeregister[17][19]~q ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hD9C8;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N11
dffeas \storeregister[29][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][19] .is_wysiwyg = "true";
defparam \storeregister[29][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N27
dffeas \storeregister[21][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][19] .is_wysiwyg = "true";
defparam \storeregister[21][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N26
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (\Mux12~0_combout  & ((\storeregister[29][19]~q ) # ((!temp_imemload_output_23)))) # (!\Mux12~0_combout  & (((\storeregister[21][19]~q  & temp_imemload_output_23))))

	.dataa(\Mux12~0_combout ),
	.datab(\storeregister[29][19]~q ),
	.datac(\storeregister[21][19]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hD8AA;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N22
cycloneive_lcell_comb \storeregister[19][19]~feeder (
// Equation(s):
// \storeregister[19][19]~feeder_combout  = Mux12

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux12),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[19][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[19][19]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[19][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N23
dffeas \storeregister[19][19] (
	.clk(!CLK),
	.d(\storeregister[19][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][19] .is_wysiwyg = "true";
defparam \storeregister[19][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N22
cycloneive_lcell_comb \storeregister[27][19]~feeder (
// Equation(s):
// \storeregister[27][19]~feeder_combout  = Mux12

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux12),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][19]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N23
dffeas \storeregister[27][19] (
	.clk(!CLK),
	.d(\storeregister[27][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][19] .is_wysiwyg = "true";
defparam \storeregister[27][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N10
cycloneive_lcell_comb \Mux12~7 (
// Equation(s):
// \Mux12~7_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[27][19]~q ))) # (!temp_imemload_output_24 & (\storeregister[19][19]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[19][19]~q ),
	.datad(\storeregister[27][19]~q ),
	.cin(gnd),
	.combout(\Mux12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~7 .lut_mask = 16'hDC98;
defparam \Mux12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N16
cycloneive_lcell_comb \storeregister[31][19]~feeder (
// Equation(s):
// \storeregister[31][19]~feeder_combout  = Mux12

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux12),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[31][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][19]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[31][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N17
dffeas \storeregister[31][19] (
	.clk(!CLK),
	.d(\storeregister[31][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][19] .is_wysiwyg = "true";
defparam \storeregister[31][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N16
cycloneive_lcell_comb \storeregister[23][19]~feeder (
// Equation(s):
// \storeregister[23][19]~feeder_combout  = Mux12

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux12),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[23][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][19]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[23][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N17
dffeas \storeregister[23][19] (
	.clk(!CLK),
	.d(\storeregister[23][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][19] .is_wysiwyg = "true";
defparam \storeregister[23][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N14
cycloneive_lcell_comb \Mux12~8 (
// Equation(s):
// \Mux12~8_combout  = (\Mux12~7_combout  & ((\storeregister[31][19]~q ) # ((!temp_imemload_output_23)))) # (!\Mux12~7_combout  & (((\storeregister[23][19]~q  & temp_imemload_output_23))))

	.dataa(\Mux12~7_combout ),
	.datab(\storeregister[31][19]~q ),
	.datac(\storeregister[23][19]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux12~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~8 .lut_mask = 16'hD8AA;
defparam \Mux12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N22
cycloneive_lcell_comb \storeregister[14][19]~feeder (
// Equation(s):
// \storeregister[14][19]~feeder_combout  = Mux12

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux12),
	.cin(gnd),
	.combout(\storeregister[14][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][19]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N23
dffeas \storeregister[14][19] (
	.clk(!CLK),
	.d(\storeregister[14][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][19] .is_wysiwyg = "true";
defparam \storeregister[14][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N28
cycloneive_lcell_comb \storeregister[15][19]~feeder (
// Equation(s):
// \storeregister[15][19]~feeder_combout  = Mux12

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux12),
	.cin(gnd),
	.combout(\storeregister[15][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][19]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N29
dffeas \storeregister[15][19] (
	.clk(!CLK),
	.d(\storeregister[15][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][19] .is_wysiwyg = "true";
defparam \storeregister[15][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N5
dffeas \storeregister[13][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][19] .is_wysiwyg = "true";
defparam \storeregister[13][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N7
dffeas \storeregister[12][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][19] .is_wysiwyg = "true";
defparam \storeregister[12][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N6
cycloneive_lcell_comb \Mux12~17 (
// Equation(s):
// \Mux12~17_combout  = (temp_imemload_output_21 & ((\storeregister[13][19]~q ) # ((temp_imemload_output_22)))) # (!temp_imemload_output_21 & (((\storeregister[12][19]~q  & !temp_imemload_output_22))))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[13][19]~q ),
	.datac(\storeregister[12][19]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux12~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~17 .lut_mask = 16'hAAD8;
defparam \Mux12~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N26
cycloneive_lcell_comb \Mux12~18 (
// Equation(s):
// \Mux12~18_combout  = (\Mux12~17_combout  & (((\storeregister[15][19]~q ) # (!temp_imemload_output_22)))) # (!\Mux12~17_combout  & (\storeregister[14][19]~q  & ((temp_imemload_output_22))))

	.dataa(\storeregister[14][19]~q ),
	.datab(\storeregister[15][19]~q ),
	.datac(\Mux12~17_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux12~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~18 .lut_mask = 16'hCAF0;
defparam \Mux12~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N25
dffeas \storeregister[9][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][19] .is_wysiwyg = "true";
defparam \storeregister[9][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N3
dffeas \storeregister[11][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][19] .is_wysiwyg = "true";
defparam \storeregister[11][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N2
cycloneive_lcell_comb \Mux12~13 (
// Equation(s):
// \Mux12~13_combout  = (\Mux12~12_combout  & (((\storeregister[11][19]~q ) # (!temp_imemload_output_21)))) # (!\Mux12~12_combout  & (\storeregister[9][19]~q  & ((temp_imemload_output_21))))

	.dataa(\Mux12~12_combout ),
	.datab(\storeregister[9][19]~q ),
	.datac(\storeregister[11][19]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux12~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~13 .lut_mask = 16'hE4AA;
defparam \Mux12~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N19
dffeas \storeregister[2][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][19] .is_wysiwyg = "true";
defparam \storeregister[2][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N19
dffeas \storeregister[1][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][19] .is_wysiwyg = "true";
defparam \storeregister[1][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N29
dffeas \storeregister[3][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][19] .is_wysiwyg = "true";
defparam \storeregister[3][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N28
cycloneive_lcell_comb \Mux12~14 (
// Equation(s):
// \Mux12~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][19]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][19]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[1][19]~q ),
	.datac(\storeregister[3][19]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux12~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~14 .lut_mask = 16'hE400;
defparam \Mux12~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N18
cycloneive_lcell_comb \Mux12~15 (
// Equation(s):
// \Mux12~15_combout  = (\Mux12~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][19]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[2][19]~q ),
	.datad(\Mux12~14_combout ),
	.cin(gnd),
	.combout(\Mux12~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~15 .lut_mask = 16'hFF40;
defparam \Mux12~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N26
cycloneive_lcell_comb \Mux12~16 (
// Equation(s):
// \Mux12~16_combout  = (temp_imemload_output_24 & ((\Mux12~13_combout ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((!temp_imemload_output_23 & \Mux12~15_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\Mux12~13_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux12~15_combout ),
	.cin(gnd),
	.combout(\Mux12~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~16 .lut_mask = 16'hADA8;
defparam \Mux12~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N22
cycloneive_lcell_comb \storeregister[6][19]~feeder (
// Equation(s):
// \storeregister[6][19]~feeder_combout  = Mux12

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux12),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[6][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[6][19]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[6][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N23
dffeas \storeregister[6][19] (
	.clk(!CLK),
	.d(\storeregister[6][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][19] .is_wysiwyg = "true";
defparam \storeregister[6][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N29
dffeas \storeregister[5][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][19] .is_wysiwyg = "true";
defparam \storeregister[5][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N28
cycloneive_lcell_comb \Mux12~10 (
// Equation(s):
// \Mux12~10_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[5][19]~q ))) # (!temp_imemload_output_21 & (\storeregister[4][19]~q ))))

	.dataa(\storeregister[4][19]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[5][19]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux12~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~10 .lut_mask = 16'hFC22;
defparam \Mux12~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N27
dffeas \storeregister[7][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][19] .is_wysiwyg = "true";
defparam \storeregister[7][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N12
cycloneive_lcell_comb \Mux12~11 (
// Equation(s):
// \Mux12~11_combout  = (\Mux12~10_combout  & (((\storeregister[7][19]~q ) # (!temp_imemload_output_22)))) # (!\Mux12~10_combout  & (\storeregister[6][19]~q  & ((temp_imemload_output_22))))

	.dataa(\storeregister[6][19]~q ),
	.datab(\Mux12~10_combout ),
	.datac(\storeregister[7][19]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux12~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~11 .lut_mask = 16'hE2CC;
defparam \Mux12~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N4
cycloneive_lcell_comb \storeregister[28][18]~feeder (
// Equation(s):
// \storeregister[28][18]~feeder_combout  = Mux13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux13),
	.cin(gnd),
	.combout(\storeregister[28][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][18]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[28][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N5
dffeas \storeregister[28][18] (
	.clk(!CLK),
	.d(\storeregister[28][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][18] .is_wysiwyg = "true";
defparam \storeregister[28][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N26
cycloneive_lcell_comb \storeregister[20][18]~feeder (
// Equation(s):
// \storeregister[20][18]~feeder_combout  = Mux13

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux13),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[20][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][18]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[20][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N27
dffeas \storeregister[20][18] (
	.clk(!CLK),
	.d(\storeregister[20][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][18] .is_wysiwyg = "true";
defparam \storeregister[20][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N17
dffeas \storeregister[24][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][18] .is_wysiwyg = "true";
defparam \storeregister[24][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N16
cycloneive_lcell_comb \Mux13~4 (
// Equation(s):
// \Mux13~4_combout  = (temp_imemload_output_24 & (((\storeregister[24][18]~q ) # (temp_imemload_output_23)))) # (!temp_imemload_output_24 & (\storeregister[16][18]~q  & ((!temp_imemload_output_23))))

	.dataa(\storeregister[16][18]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[24][18]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~4 .lut_mask = 16'hCCE2;
defparam \Mux13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N26
cycloneive_lcell_comb \Mux13~5 (
// Equation(s):
// \Mux13~5_combout  = (temp_imemload_output_23 & ((\Mux13~4_combout  & (\storeregister[28][18]~q )) # (!\Mux13~4_combout  & ((\storeregister[20][18]~q ))))) # (!temp_imemload_output_23 & (((\Mux13~4_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[28][18]~q ),
	.datac(\storeregister[20][18]~q ),
	.datad(\Mux13~4_combout ),
	.cin(gnd),
	.combout(\Mux13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~5 .lut_mask = 16'hDDA0;
defparam \Mux13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N9
dffeas \storeregister[30][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][18] .is_wysiwyg = "true";
defparam \storeregister[30][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N6
cycloneive_lcell_comb \storeregister[22][18]~feeder (
// Equation(s):
// \storeregister[22][18]~feeder_combout  = Mux13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux13),
	.cin(gnd),
	.combout(\storeregister[22][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[22][18]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[22][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N7
dffeas \storeregister[22][18] (
	.clk(!CLK),
	.d(\storeregister[22][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][18] .is_wysiwyg = "true";
defparam \storeregister[22][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N8
cycloneive_lcell_comb \Mux13~3 (
// Equation(s):
// \Mux13~3_combout  = (\Mux13~2_combout  & (((\storeregister[30][18]~q )) # (!temp_imemload_output_23))) # (!\Mux13~2_combout  & (temp_imemload_output_23 & ((\storeregister[22][18]~q ))))

	.dataa(\Mux13~2_combout ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[30][18]~q ),
	.datad(\storeregister[22][18]~q ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~3 .lut_mask = 16'hE6A2;
defparam \Mux13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N12
cycloneive_lcell_comb \Mux13~6 (
// Equation(s):
// \Mux13~6_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & ((\Mux13~3_combout ))) # (!temp_imemload_output_22 & (\Mux13~5_combout ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\Mux13~5_combout ),
	.datad(\Mux13~3_combout ),
	.cin(gnd),
	.combout(\Mux13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~6 .lut_mask = 16'hDC98;
defparam \Mux13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N31
dffeas \storeregister[27][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][18] .is_wysiwyg = "true";
defparam \storeregister[27][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N29
dffeas \storeregister[31][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][18] .is_wysiwyg = "true";
defparam \storeregister[31][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N17
dffeas \storeregister[23][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][18] .is_wysiwyg = "true";
defparam \storeregister[23][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N19
dffeas \storeregister[19][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][18] .is_wysiwyg = "true";
defparam \storeregister[19][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N18
cycloneive_lcell_comb \Mux13~7 (
// Equation(s):
// \Mux13~7_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[23][18]~q )) # (!temp_imemload_output_23 & ((\storeregister[19][18]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[23][18]~q ),
	.datac(\storeregister[19][18]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~7 .lut_mask = 16'hEE50;
defparam \Mux13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N28
cycloneive_lcell_comb \Mux13~8 (
// Equation(s):
// \Mux13~8_combout  = (temp_imemload_output_24 & ((\Mux13~7_combout  & ((\storeregister[31][18]~q ))) # (!\Mux13~7_combout  & (\storeregister[27][18]~q )))) # (!temp_imemload_output_24 & (((\Mux13~7_combout ))))

	.dataa(\storeregister[27][18]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[31][18]~q ),
	.datad(\Mux13~7_combout ),
	.cin(gnd),
	.combout(\Mux13~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~8 .lut_mask = 16'hF388;
defparam \Mux13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N23
dffeas \storeregister[29][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][18] .is_wysiwyg = "true";
defparam \storeregister[29][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N24
cycloneive_lcell_comb \storeregister[17][18]~feeder (
// Equation(s):
// \storeregister[17][18]~feeder_combout  = Mux13

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux13),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[17][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[17][18]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[17][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N25
dffeas \storeregister[17][18] (
	.clk(!CLK),
	.d(\storeregister[17][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][18] .is_wysiwyg = "true";
defparam \storeregister[17][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N25
dffeas \storeregister[21][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][18] .is_wysiwyg = "true";
defparam \storeregister[21][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N24
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[21][18]~q ))) # (!temp_imemload_output_23 & (\storeregister[17][18]~q ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[17][18]~q ),
	.datac(\storeregister[21][18]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hFA44;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N21
dffeas \storeregister[25][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][18] .is_wysiwyg = "true";
defparam \storeregister[25][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N20
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (\Mux13~0_combout  & ((\storeregister[29][18]~q ) # ((!temp_imemload_output_24)))) # (!\Mux13~0_combout  & (((\storeregister[25][18]~q  & temp_imemload_output_24))))

	.dataa(\storeregister[29][18]~q ),
	.datab(\Mux13~0_combout ),
	.datac(\storeregister[25][18]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hB8CC;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N10
cycloneive_lcell_comb \storeregister[15][18]~feeder (
// Equation(s):
// \storeregister[15][18]~feeder_combout  = Mux13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux13),
	.cin(gnd),
	.combout(\storeregister[15][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][18]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N11
dffeas \storeregister[15][18] (
	.clk(!CLK),
	.d(\storeregister[15][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][18] .is_wysiwyg = "true";
defparam \storeregister[15][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N20
cycloneive_lcell_comb \storeregister[14][18]~feeder (
// Equation(s):
// \storeregister[14][18]~feeder_combout  = Mux13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux13),
	.cin(gnd),
	.combout(\storeregister[14][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][18]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y40_N21
dffeas \storeregister[14][18] (
	.clk(!CLK),
	.d(\storeregister[14][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][18] .is_wysiwyg = "true";
defparam \storeregister[14][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N25
dffeas \storeregister[13][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][18] .is_wysiwyg = "true";
defparam \storeregister[13][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N11
dffeas \storeregister[12][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][18] .is_wysiwyg = "true";
defparam \storeregister[12][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N24
cycloneive_lcell_comb \Mux13~17 (
// Equation(s):
// \Mux13~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][18]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[12][18]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[13][18]~q ),
	.datad(\storeregister[12][18]~q ),
	.cin(gnd),
	.combout(\Mux13~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~17 .lut_mask = 16'hB9A8;
defparam \Mux13~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N8
cycloneive_lcell_comb \Mux13~18 (
// Equation(s):
// \Mux13~18_combout  = (temp_imemload_output_22 & ((\Mux13~17_combout  & (\storeregister[15][18]~q )) # (!\Mux13~17_combout  & ((\storeregister[14][18]~q ))))) # (!temp_imemload_output_22 & (((\Mux13~17_combout ))))

	.dataa(\storeregister[15][18]~q ),
	.datab(\storeregister[14][18]~q ),
	.datac(temp_imemload_output_22),
	.datad(\Mux13~17_combout ),
	.cin(gnd),
	.combout(\Mux13~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~18 .lut_mask = 16'hAFC0;
defparam \Mux13~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N23
dffeas \storeregister[11][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][18] .is_wysiwyg = "true";
defparam \storeregister[11][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N19
dffeas \storeregister[10][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][18] .is_wysiwyg = "true";
defparam \storeregister[10][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N13
dffeas \storeregister[8][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][18] .is_wysiwyg = "true";
defparam \storeregister[8][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N18
cycloneive_lcell_comb \Mux13~10 (
// Equation(s):
// \Mux13~10_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\storeregister[10][18]~q )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & ((\storeregister[8][18]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[10][18]~q ),
	.datad(\storeregister[8][18]~q ),
	.cin(gnd),
	.combout(\Mux13~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~10 .lut_mask = 16'hB9A8;
defparam \Mux13~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N17
dffeas \storeregister[9][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][18] .is_wysiwyg = "true";
defparam \storeregister[9][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N16
cycloneive_lcell_comb \Mux13~11 (
// Equation(s):
// \Mux13~11_combout  = (\Mux13~10_combout  & ((\storeregister[11][18]~q ) # ((!temp_imemload_output_21)))) # (!\Mux13~10_combout  & (((\storeregister[9][18]~q  & temp_imemload_output_21))))

	.dataa(\storeregister[11][18]~q ),
	.datab(\Mux13~10_combout ),
	.datac(\storeregister[9][18]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux13~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~11 .lut_mask = 16'hB8CC;
defparam \Mux13~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N18
cycloneive_lcell_comb \storeregister[2][18]~feeder (
// Equation(s):
// \storeregister[2][18]~feeder_combout  = Mux13

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux13),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[2][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[2][18]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[2][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N19
dffeas \storeregister[2][18] (
	.clk(!CLK),
	.d(\storeregister[2][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][18] .is_wysiwyg = "true";
defparam \storeregister[2][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N8
cycloneive_lcell_comb \Mux13~15 (
// Equation(s):
// \Mux13~15_combout  = (\Mux13~14_combout ) # ((\storeregister[2][18]~q  & (!temp_imemload_output_21 & temp_imemload_output_22)))

	.dataa(\Mux13~14_combout ),
	.datab(\storeregister[2][18]~q ),
	.datac(temp_imemload_output_21),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux13~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~15 .lut_mask = 16'hAEAA;
defparam \Mux13~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y40_N11
dffeas \storeregister[4][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][18] .is_wysiwyg = "true";
defparam \storeregister[4][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y40_N1
dffeas \storeregister[5][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][18] .is_wysiwyg = "true";
defparam \storeregister[5][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N10
cycloneive_lcell_comb \Mux13~12 (
// Equation(s):
// \Mux13~12_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[5][18]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & (\storeregister[4][18]~q )))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[4][18]~q ),
	.datad(\storeregister[5][18]~q ),
	.cin(gnd),
	.combout(\Mux13~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~12 .lut_mask = 16'hBA98;
defparam \Mux13~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N21
dffeas \storeregister[7][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][18] .is_wysiwyg = "true";
defparam \storeregister[7][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N11
dffeas \storeregister[6][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][18] .is_wysiwyg = "true";
defparam \storeregister[6][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N20
cycloneive_lcell_comb \Mux13~13 (
// Equation(s):
// \Mux13~13_combout  = (temp_imemload_output_22 & ((\Mux13~12_combout  & (\storeregister[7][18]~q )) # (!\Mux13~12_combout  & ((\storeregister[6][18]~q ))))) # (!temp_imemload_output_22 & (\Mux13~12_combout ))

	.dataa(temp_imemload_output_22),
	.datab(\Mux13~12_combout ),
	.datac(\storeregister[7][18]~q ),
	.datad(\storeregister[6][18]~q ),
	.cin(gnd),
	.combout(\Mux13~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~13 .lut_mask = 16'hE6C4;
defparam \Mux13~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N0
cycloneive_lcell_comb \Mux13~16 (
// Equation(s):
// \Mux13~16_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\Mux13~13_combout ))) # (!temp_imemload_output_23 & (\Mux13~15_combout ))))

	.dataa(\Mux13~15_combout ),
	.datab(temp_imemload_output_24),
	.datac(\Mux13~13_combout ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux13~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~16 .lut_mask = 16'hFC22;
defparam \Mux13~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N1
dffeas \storeregister[29][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][24] .is_wysiwyg = "true";
defparam \storeregister[29][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N13
dffeas \storeregister[25][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][24] .is_wysiwyg = "true";
defparam \storeregister[25][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N19
dffeas \storeregister[21][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][24] .is_wysiwyg = "true";
defparam \storeregister[21][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N18
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[21][24]~q ))) # (!temp_imemload_output_23 & (\storeregister[17][24]~q ))))

	.dataa(\storeregister[17][24]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[21][24]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hFC22;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N12
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (temp_imemload_output_24 & ((\Mux7~0_combout  & (\storeregister[29][24]~q )) # (!\Mux7~0_combout  & ((\storeregister[25][24]~q ))))) # (!temp_imemload_output_24 & (((\Mux7~0_combout ))))

	.dataa(\storeregister[29][24]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[25][24]~q ),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hBBC0;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N19
dffeas \storeregister[19][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][24] .is_wysiwyg = "true";
defparam \storeregister[19][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N18
cycloneive_lcell_comb \Mux7~7 (
// Equation(s):
// \Mux7~7_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[23][24]~q )) # (!temp_imemload_output_23 & ((\storeregister[19][24]~q )))))

	.dataa(\storeregister[23][24]~q ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[19][24]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~7 .lut_mask = 16'hEE30;
defparam \Mux7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N16
cycloneive_lcell_comb \storeregister[31][24]~feeder (
// Equation(s):
// \storeregister[31][24]~feeder_combout  = Mux7

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux7),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[31][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[31][24]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[31][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N17
dffeas \storeregister[31][24] (
	.clk(!CLK),
	.d(\storeregister[31][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][24] .is_wysiwyg = "true";
defparam \storeregister[31][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N25
dffeas \storeregister[27][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][24] .is_wysiwyg = "true";
defparam \storeregister[27][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N30
cycloneive_lcell_comb \Mux7~8 (
// Equation(s):
// \Mux7~8_combout  = (\Mux7~7_combout  & ((\storeregister[31][24]~q ) # ((!temp_imemload_output_24)))) # (!\Mux7~7_combout  & (((\storeregister[27][24]~q  & temp_imemload_output_24))))

	.dataa(\Mux7~7_combout ),
	.datab(\storeregister[31][24]~q ),
	.datac(\storeregister[27][24]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~8 .lut_mask = 16'hD8AA;
defparam \Mux7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N24
cycloneive_lcell_comb \storeregister[30][24]~feeder (
// Equation(s):
// \storeregister[30][24]~feeder_combout  = Mux7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux7),
	.cin(gnd),
	.combout(\storeregister[30][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[30][24]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[30][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N25
dffeas \storeregister[30][24] (
	.clk(!CLK),
	.d(\storeregister[30][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][24] .is_wysiwyg = "true";
defparam \storeregister[30][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N9
dffeas \storeregister[26][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][24] .is_wysiwyg = "true";
defparam \storeregister[26][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N19
dffeas \storeregister[18][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][24] .is_wysiwyg = "true";
defparam \storeregister[18][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N18
cycloneive_lcell_comb \Mux7~2 (
// Equation(s):
// \Mux7~2_combout  = (temp_imemload_output_24 & ((\storeregister[26][24]~q ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((\storeregister[18][24]~q  & !temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[26][24]~q ),
	.datac(\storeregister[18][24]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~2 .lut_mask = 16'hAAD8;
defparam \Mux7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N30
cycloneive_lcell_comb \Mux7~3 (
// Equation(s):
// \Mux7~3_combout  = (temp_imemload_output_23 & ((\Mux7~2_combout  & ((\storeregister[30][24]~q ))) # (!\Mux7~2_combout  & (\storeregister[22][24]~q )))) # (!temp_imemload_output_23 & (((\Mux7~2_combout ))))

	.dataa(\storeregister[22][24]~q ),
	.datab(\storeregister[30][24]~q ),
	.datac(temp_imemload_output_23),
	.datad(\Mux7~2_combout ),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~3 .lut_mask = 16'hCFA0;
defparam \Mux7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N22
cycloneive_lcell_comb \storeregister[28][24]~feeder (
// Equation(s):
// \storeregister[28][24]~feeder_combout  = Mux7

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux7),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[28][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][24]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[28][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N23
dffeas \storeregister[28][24] (
	.clk(!CLK),
	.d(\storeregister[28][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][24] .is_wysiwyg = "true";
defparam \storeregister[28][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N15
dffeas \storeregister[16][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][24] .is_wysiwyg = "true";
defparam \storeregister[16][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N20
cycloneive_lcell_comb \storeregister[24][24]~feeder (
// Equation(s):
// \storeregister[24][24]~feeder_combout  = Mux7

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux7),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[24][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][24]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[24][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N21
dffeas \storeregister[24][24] (
	.clk(!CLK),
	.d(\storeregister[24][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][24] .is_wysiwyg = "true";
defparam \storeregister[24][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N24
cycloneive_lcell_comb \Mux7~4 (
// Equation(s):
// \Mux7~4_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[24][24]~q ))) # (!temp_imemload_output_24 & (\storeregister[16][24]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][24]~q ),
	.datad(\storeregister[24][24]~q ),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~4 .lut_mask = 16'hDC98;
defparam \Mux7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N22
cycloneive_lcell_comb \Mux7~5 (
// Equation(s):
// \Mux7~5_combout  = (temp_imemload_output_23 & ((\Mux7~4_combout  & ((\storeregister[28][24]~q ))) # (!\Mux7~4_combout  & (\storeregister[20][24]~q )))) # (!temp_imemload_output_23 & (((\Mux7~4_combout ))))

	.dataa(\storeregister[20][24]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[28][24]~q ),
	.datad(\Mux7~4_combout ),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~5 .lut_mask = 16'hF388;
defparam \Mux7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N16
cycloneive_lcell_comb \Mux7~6 (
// Equation(s):
// \Mux7~6_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\Mux7~3_combout )) # (!temp_imemload_output_22 & ((\Mux7~5_combout )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\Mux7~3_combout ),
	.datad(\Mux7~5_combout ),
	.cin(gnd),
	.combout(\Mux7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~6 .lut_mask = 16'hD9C8;
defparam \Mux7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N5
dffeas \storeregister[13][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][24] .is_wysiwyg = "true";
defparam \storeregister[13][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N4
cycloneive_lcell_comb \Mux7~17 (
// Equation(s):
// \Mux7~17_combout  = (temp_imemload_output_22 & (((temp_imemload_output_21)))) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[13][24]~q ))) # (!temp_imemload_output_21 & (\storeregister[12][24]~q ))))

	.dataa(\storeregister[12][24]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[13][24]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux7~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~17 .lut_mask = 16'hFC22;
defparam \Mux7~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N4
cycloneive_lcell_comb \storeregister[14][24]~feeder (
// Equation(s):
// \storeregister[14][24]~feeder_combout  = Mux7

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux7),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[14][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][24]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[14][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y43_N5
dffeas \storeregister[14][24] (
	.clk(!CLK),
	.d(\storeregister[14][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][24] .is_wysiwyg = "true";
defparam \storeregister[14][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N2
cycloneive_lcell_comb \storeregister[15][24]~feeder (
// Equation(s):
// \storeregister[15][24]~feeder_combout  = Mux7

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux7),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[15][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][24]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[15][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y43_N3
dffeas \storeregister[15][24] (
	.clk(!CLK),
	.d(\storeregister[15][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][24] .is_wysiwyg = "true";
defparam \storeregister[15][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N8
cycloneive_lcell_comb \Mux7~18 (
// Equation(s):
// \Mux7~18_combout  = (\Mux7~17_combout  & (((\storeregister[15][24]~q ) # (!temp_imemload_output_22)))) # (!\Mux7~17_combout  & (\storeregister[14][24]~q  & (temp_imemload_output_22)))

	.dataa(\Mux7~17_combout ),
	.datab(\storeregister[14][24]~q ),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[15][24]~q ),
	.cin(gnd),
	.combout(\Mux7~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~18 .lut_mask = 16'hEA4A;
defparam \Mux7~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N21
dffeas \storeregister[10][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][24] .is_wysiwyg = "true";
defparam \storeregister[10][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N21
dffeas \storeregister[8][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][24] .is_wysiwyg = "true";
defparam \storeregister[8][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N20
cycloneive_lcell_comb \Mux7~10 (
// Equation(s):
// \Mux7~10_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[10][24]~q )) # (!temp_imemload_output_22 & ((\storeregister[8][24]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][24]~q ),
	.datad(\storeregister[8][24]~q ),
	.cin(gnd),
	.combout(\Mux7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~10 .lut_mask = 16'hD9C8;
defparam \Mux7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N23
dffeas \storeregister[9][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][24] .is_wysiwyg = "true";
defparam \storeregister[9][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N31
dffeas \storeregister[11][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][24] .is_wysiwyg = "true";
defparam \storeregister[11][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N22
cycloneive_lcell_comb \Mux7~11 (
// Equation(s):
// \Mux7~11_combout  = (\Mux7~10_combout  & (((\storeregister[11][24]~q )) # (!temp_imemload_output_21))) # (!\Mux7~10_combout  & (temp_imemload_output_21 & (\storeregister[9][24]~q )))

	.dataa(\Mux7~10_combout ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[9][24]~q ),
	.datad(\storeregister[11][24]~q ),
	.cin(gnd),
	.combout(\Mux7~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~11 .lut_mask = 16'hEA62;
defparam \Mux7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y41_N15
dffeas \storeregister[4][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][24] .is_wysiwyg = "true";
defparam \storeregister[4][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N14
cycloneive_lcell_comb \Mux7~12 (
// Equation(s):
// \Mux7~12_combout  = (temp_imemload_output_21 & ((\storeregister[5][24]~q ) # ((temp_imemload_output_22)))) # (!temp_imemload_output_21 & (((\storeregister[4][24]~q  & !temp_imemload_output_22))))

	.dataa(\storeregister[5][24]~q ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[4][24]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux7~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~12 .lut_mask = 16'hCCB8;
defparam \Mux7~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N9
dffeas \storeregister[7][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][24] .is_wysiwyg = "true";
defparam \storeregister[7][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N8
cycloneive_lcell_comb \Mux7~13 (
// Equation(s):
// \Mux7~13_combout  = (\Mux7~12_combout  & (((\storeregister[7][24]~q ) # (!temp_imemload_output_22)))) # (!\Mux7~12_combout  & (\storeregister[6][24]~q  & ((temp_imemload_output_22))))

	.dataa(\storeregister[6][24]~q ),
	.datab(\Mux7~12_combout ),
	.datac(\storeregister[7][24]~q ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux7~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~13 .lut_mask = 16'hE2CC;
defparam \Mux7~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N26
cycloneive_lcell_comb \storeregister[2][24]~feeder (
// Equation(s):
// \storeregister[2][24]~feeder_combout  = Mux7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux7),
	.cin(gnd),
	.combout(\storeregister[2][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[2][24]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[2][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y42_N27
dffeas \storeregister[2][24] (
	.clk(!CLK),
	.d(\storeregister[2][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][24] .is_wysiwyg = "true";
defparam \storeregister[2][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N29
dffeas \storeregister[3][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][24] .is_wysiwyg = "true";
defparam \storeregister[3][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N28
cycloneive_lcell_comb \Mux7~14 (
// Equation(s):
// \Mux7~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & ((\storeregister[3][24]~q ))) # (!temp_imemload_output_22 & (\storeregister[1][24]~q ))))

	.dataa(\storeregister[1][24]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[3][24]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux7~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~14 .lut_mask = 16'hE200;
defparam \Mux7~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N8
cycloneive_lcell_comb \Mux7~15 (
// Equation(s):
// \Mux7~15_combout  = (\Mux7~14_combout ) # ((temp_imemload_output_22 & (!temp_imemload_output_21 & \storeregister[2][24]~q )))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[2][24]~q ),
	.datad(\Mux7~14_combout ),
	.cin(gnd),
	.combout(\Mux7~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~15 .lut_mask = 16'hFF20;
defparam \Mux7~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N16
cycloneive_lcell_comb \Mux7~16 (
// Equation(s):
// \Mux7~16_combout  = (temp_imemload_output_23 & ((\Mux7~13_combout ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\Mux7~15_combout  & !temp_imemload_output_24))))

	.dataa(\Mux7~13_combout ),
	.datab(temp_imemload_output_23),
	.datac(\Mux7~15_combout ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux7~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~16 .lut_mask = 16'hCCB8;
defparam \Mux7~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N7
dffeas \storeregister[30][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][23] .is_wysiwyg = "true";
defparam \storeregister[30][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N29
dffeas \storeregister[26][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][23] .is_wysiwyg = "true";
defparam \storeregister[26][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N6
cycloneive_lcell_comb \Mux8~3 (
// Equation(s):
// \Mux8~3_combout  = (\Mux8~2_combout  & (((\storeregister[30][23]~q )) # (!temp_imemload_output_24))) # (!\Mux8~2_combout  & (temp_imemload_output_24 & ((\storeregister[26][23]~q ))))

	.dataa(\Mux8~2_combout ),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[30][23]~q ),
	.datad(\storeregister[26][23]~q ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~3 .lut_mask = 16'hE6A2;
defparam \Mux8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N28
cycloneive_lcell_comb \storeregister[28][23]~feeder (
// Equation(s):
// \storeregister[28][23]~feeder_combout  = Mux8

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux8),
	.cin(gnd),
	.combout(\storeregister[28][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][23]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[28][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N29
dffeas \storeregister[28][23] (
	.clk(!CLK),
	.d(\storeregister[28][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][23] .is_wysiwyg = "true";
defparam \storeregister[28][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N9
dffeas \storeregister[24][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][23] .is_wysiwyg = "true";
defparam \storeregister[24][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N27
dffeas \storeregister[16][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][23] .is_wysiwyg = "true";
defparam \storeregister[16][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N21
dffeas \storeregister[20][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][23] .is_wysiwyg = "true";
defparam \storeregister[20][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N26
cycloneive_lcell_comb \Mux8~4 (
// Equation(s):
// \Mux8~4_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & ((\storeregister[20][23]~q ))) # (!temp_imemload_output_23 & (\storeregister[16][23]~q ))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[16][23]~q ),
	.datad(\storeregister[20][23]~q ),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~4 .lut_mask = 16'hDC98;
defparam \Mux8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N10
cycloneive_lcell_comb \Mux8~5 (
// Equation(s):
// \Mux8~5_combout  = (temp_imemload_output_24 & ((\Mux8~4_combout  & (\storeregister[28][23]~q )) # (!\Mux8~4_combout  & ((\storeregister[24][23]~q ))))) # (!temp_imemload_output_24 & (((\Mux8~4_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[28][23]~q ),
	.datac(\storeregister[24][23]~q ),
	.datad(\Mux8~4_combout ),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~5 .lut_mask = 16'hDDA0;
defparam \Mux8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N30
cycloneive_lcell_comb \Mux8~6 (
// Equation(s):
// \Mux8~6_combout  = (temp_imemload_output_21 & (temp_imemload_output_22)) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & (\Mux8~3_combout )) # (!temp_imemload_output_22 & ((\Mux8~5_combout )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\Mux8~3_combout ),
	.datad(\Mux8~5_combout ),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~6 .lut_mask = 16'hD9C8;
defparam \Mux8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N20
cycloneive_lcell_comb \storeregister[21][23]~feeder (
// Equation(s):
// \storeregister[21][23]~feeder_combout  = Mux8

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux8),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[21][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][23]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[21][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N21
dffeas \storeregister[21][23] (
	.clk(!CLK),
	.d(\storeregister[21][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][23] .is_wysiwyg = "true";
defparam \storeregister[21][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N19
dffeas \storeregister[29][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][23] .is_wysiwyg = "true";
defparam \storeregister[29][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N5
dffeas \storeregister[25][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][23] .is_wysiwyg = "true";
defparam \storeregister[25][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N17
dffeas \storeregister[17][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][23] .is_wysiwyg = "true";
defparam \storeregister[17][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N16
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[25][23]~q )) # (!temp_imemload_output_24 & ((\storeregister[17][23]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[25][23]~q ),
	.datac(\storeregister[17][23]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hEE50;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N18
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (temp_imemload_output_23 & ((\Mux8~0_combout  & ((\storeregister[29][23]~q ))) # (!\Mux8~0_combout  & (\storeregister[21][23]~q )))) # (!temp_imemload_output_23 & (((\Mux8~0_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[21][23]~q ),
	.datac(\storeregister[29][23]~q ),
	.datad(\Mux8~0_combout ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hF588;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N29
dffeas \storeregister[23][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][23] .is_wysiwyg = "true";
defparam \storeregister[23][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N10
cycloneive_lcell_comb \storeregister[19][23]~feeder (
// Equation(s):
// \storeregister[19][23]~feeder_combout  = Mux8

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux8),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[19][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[19][23]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[19][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N11
dffeas \storeregister[19][23] (
	.clk(!CLK),
	.d(\storeregister[19][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][23] .is_wysiwyg = "true";
defparam \storeregister[19][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N23
dffeas \storeregister[27][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][23] .is_wysiwyg = "true";
defparam \storeregister[27][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N22
cycloneive_lcell_comb \Mux8~7 (
// Equation(s):
// \Mux8~7_combout  = (temp_imemload_output_24 & (((\storeregister[27][23]~q ) # (temp_imemload_output_23)))) # (!temp_imemload_output_24 & (\storeregister[19][23]~q  & ((!temp_imemload_output_23))))

	.dataa(temp_imemload_output_24),
	.datab(\storeregister[19][23]~q ),
	.datac(\storeregister[27][23]~q ),
	.datad(temp_imemload_output_23),
	.cin(gnd),
	.combout(\Mux8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~7 .lut_mask = 16'hAAE4;
defparam \Mux8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N17
dffeas \storeregister[31][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][23] .is_wysiwyg = "true";
defparam \storeregister[31][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N30
cycloneive_lcell_comb \Mux8~8 (
// Equation(s):
// \Mux8~8_combout  = (temp_imemload_output_23 & ((\Mux8~7_combout  & ((\storeregister[31][23]~q ))) # (!\Mux8~7_combout  & (\storeregister[23][23]~q )))) # (!temp_imemload_output_23 & (((\Mux8~7_combout ))))

	.dataa(\storeregister[23][23]~q ),
	.datab(temp_imemload_output_23),
	.datac(\Mux8~7_combout ),
	.datad(\storeregister[31][23]~q ),
	.cin(gnd),
	.combout(\Mux8~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~8 .lut_mask = 16'hF838;
defparam \Mux8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y41_N17
dffeas \storeregister[5][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][23] .is_wysiwyg = "true";
defparam \storeregister[5][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y41_N11
dffeas \storeregister[4][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][23] .is_wysiwyg = "true";
defparam \storeregister[4][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N16
cycloneive_lcell_comb \Mux8~10 (
// Equation(s):
// \Mux8~10_combout  = (temp_imemload_output_22 & (temp_imemload_output_21)) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & (\storeregister[5][23]~q )) # (!temp_imemload_output_21 & ((\storeregister[4][23]~q )))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[5][23]~q ),
	.datad(\storeregister[4][23]~q ),
	.cin(gnd),
	.combout(\Mux8~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~10 .lut_mask = 16'hD9C8;
defparam \Mux8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y40_N17
dffeas \storeregister[6][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][23] .is_wysiwyg = "true";
defparam \storeregister[6][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y40_N15
dffeas \storeregister[7][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][23] .is_wysiwyg = "true";
defparam \storeregister[7][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N16
cycloneive_lcell_comb \Mux8~11 (
// Equation(s):
// \Mux8~11_combout  = (\Mux8~10_combout  & (((\storeregister[7][23]~q )) # (!temp_imemload_output_22))) # (!\Mux8~10_combout  & (temp_imemload_output_22 & (\storeregister[6][23]~q )))

	.dataa(\Mux8~10_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[6][23]~q ),
	.datad(\storeregister[7][23]~q ),
	.cin(gnd),
	.combout(\Mux8~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~11 .lut_mask = 16'hEA62;
defparam \Mux8~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N12
cycloneive_lcell_comb \storeregister[2][23]~feeder (
// Equation(s):
// \storeregister[2][23]~feeder_combout  = Mux8

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux8),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[2][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[2][23]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[2][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N13
dffeas \storeregister[2][23] (
	.clk(!CLK),
	.d(\storeregister[2][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][23] .is_wysiwyg = "true";
defparam \storeregister[2][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N5
dffeas \storeregister[3][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][23] .is_wysiwyg = "true";
defparam \storeregister[3][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N19
dffeas \storeregister[1][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][23] .is_wysiwyg = "true";
defparam \storeregister[1][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N4
cycloneive_lcell_comb \Mux8~14 (
// Equation(s):
// \Mux8~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[3][23]~q )) # (!temp_imemload_output_22 & ((\storeregister[1][23]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[3][23]~q ),
	.datad(\storeregister[1][23]~q ),
	.cin(gnd),
	.combout(\Mux8~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~14 .lut_mask = 16'hA280;
defparam \Mux8~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N26
cycloneive_lcell_comb \Mux8~15 (
// Equation(s):
// \Mux8~15_combout  = (\Mux8~14_combout ) # ((!temp_imemload_output_21 & (\storeregister[2][23]~q  & temp_imemload_output_22)))

	.dataa(temp_imemload_output_21),
	.datab(\storeregister[2][23]~q ),
	.datac(\Mux8~14_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux8~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~15 .lut_mask = 16'hF4F0;
defparam \Mux8~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N15
dffeas \storeregister[11][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][23] .is_wysiwyg = "true";
defparam \storeregister[11][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N21
dffeas \storeregister[9][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][23] .is_wysiwyg = "true";
defparam \storeregister[9][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N14
cycloneive_lcell_comb \Mux8~13 (
// Equation(s):
// \Mux8~13_combout  = (\Mux8~12_combout  & (((\storeregister[11][23]~q )) # (!temp_imemload_output_21))) # (!\Mux8~12_combout  & (temp_imemload_output_21 & ((\storeregister[9][23]~q ))))

	.dataa(\Mux8~12_combout ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[11][23]~q ),
	.datad(\storeregister[9][23]~q ),
	.cin(gnd),
	.combout(\Mux8~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~13 .lut_mask = 16'hE6A2;
defparam \Mux8~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N8
cycloneive_lcell_comb \Mux8~16 (
// Equation(s):
// \Mux8~16_combout  = (temp_imemload_output_24 & ((temp_imemload_output_23) # ((\Mux8~13_combout )))) # (!temp_imemload_output_24 & (!temp_imemload_output_23 & (\Mux8~15_combout )))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\Mux8~15_combout ),
	.datad(\Mux8~13_combout ),
	.cin(gnd),
	.combout(\Mux8~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~16 .lut_mask = 16'hBA98;
defparam \Mux8~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N29
dffeas \storeregister[13][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][23] .is_wysiwyg = "true";
defparam \storeregister[13][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N7
dffeas \storeregister[12][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][23] .is_wysiwyg = "true";
defparam \storeregister[12][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N28
cycloneive_lcell_comb \Mux8~17 (
// Equation(s):
// \Mux8~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][23]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[12][23]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[13][23]~q ),
	.datad(\storeregister[12][23]~q ),
	.cin(gnd),
	.combout(\Mux8~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~17 .lut_mask = 16'hB9A8;
defparam \Mux8~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N22
cycloneive_lcell_comb \storeregister[14][23]~feeder (
// Equation(s):
// \storeregister[14][23]~feeder_combout  = Mux8

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux8),
	.cin(gnd),
	.combout(\storeregister[14][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][23]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N23
dffeas \storeregister[14][23] (
	.clk(!CLK),
	.d(\storeregister[14][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][23] .is_wysiwyg = "true";
defparam \storeregister[14][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N20
cycloneive_lcell_comb \storeregister[15][23]~feeder (
// Equation(s):
// \storeregister[15][23]~feeder_combout  = Mux8

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux8),
	.cin(gnd),
	.combout(\storeregister[15][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][23]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[15][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N21
dffeas \storeregister[15][23] (
	.clk(!CLK),
	.d(\storeregister[15][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][23] .is_wysiwyg = "true";
defparam \storeregister[15][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N2
cycloneive_lcell_comb \Mux8~18 (
// Equation(s):
// \Mux8~18_combout  = (\Mux8~17_combout  & (((\storeregister[15][23]~q )) # (!temp_imemload_output_22))) # (!\Mux8~17_combout  & (temp_imemload_output_22 & (\storeregister[14][23]~q )))

	.dataa(\Mux8~17_combout ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[14][23]~q ),
	.datad(\storeregister[15][23]~q ),
	.cin(gnd),
	.combout(\Mux8~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~18 .lut_mask = 16'hEA62;
defparam \Mux8~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N13
dffeas \storeregister[27][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][22] .is_wysiwyg = "true";
defparam \storeregister[27][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N23
dffeas \storeregister[19][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][22] .is_wysiwyg = "true";
defparam \storeregister[19][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N0
cycloneive_lcell_comb \storeregister[23][22]~feeder (
// Equation(s):
// \storeregister[23][22]~feeder_combout  = Mux9

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux9),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[23][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][22]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[23][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N1
dffeas \storeregister[23][22] (
	.clk(!CLK),
	.d(\storeregister[23][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][22] .is_wysiwyg = "true";
defparam \storeregister[23][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N22
cycloneive_lcell_comb \Mux9~7 (
// Equation(s):
// \Mux9~7_combout  = (temp_imemload_output_23 & ((temp_imemload_output_24) # ((\storeregister[23][22]~q )))) # (!temp_imemload_output_23 & (!temp_imemload_output_24 & (\storeregister[19][22]~q )))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[19][22]~q ),
	.datad(\storeregister[23][22]~q ),
	.cin(gnd),
	.combout(\Mux9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~7 .lut_mask = 16'hBA98;
defparam \Mux9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N1
dffeas \storeregister[31][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][22] .is_wysiwyg = "true";
defparam \storeregister[31][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N30
cycloneive_lcell_comb \Mux9~8 (
// Equation(s):
// \Mux9~8_combout  = (\Mux9~7_combout  & (((\storeregister[31][22]~q ) # (!temp_imemload_output_24)))) # (!\Mux9~7_combout  & (\storeregister[27][22]~q  & (temp_imemload_output_24)))

	.dataa(\storeregister[27][22]~q ),
	.datab(\Mux9~7_combout ),
	.datac(temp_imemload_output_24),
	.datad(\storeregister[31][22]~q ),
	.cin(gnd),
	.combout(\Mux9~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~8 .lut_mask = 16'hEC2C;
defparam \Mux9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N27
dffeas \storeregister[25][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][22] .is_wysiwyg = "true";
defparam \storeregister[25][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N3
dffeas \storeregister[17][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][22] .is_wysiwyg = "true";
defparam \storeregister[17][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N2
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (temp_imemload_output_23 & ((\storeregister[21][22]~q ) # ((temp_imemload_output_24)))) # (!temp_imemload_output_23 & (((\storeregister[17][22]~q  & !temp_imemload_output_24))))

	.dataa(\storeregister[21][22]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[17][22]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hCCB8;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N17
dffeas \storeregister[29][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][22] .is_wysiwyg = "true";
defparam \storeregister[29][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N16
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (\Mux9~0_combout  & (((\storeregister[29][22]~q ) # (!temp_imemload_output_24)))) # (!\Mux9~0_combout  & (\storeregister[25][22]~q  & ((temp_imemload_output_24))))

	.dataa(\storeregister[25][22]~q ),
	.datab(\Mux9~0_combout ),
	.datac(\storeregister[29][22]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hE2CC;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N31
dffeas \storeregister[30][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][22] .is_wysiwyg = "true";
defparam \storeregister[30][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N25
dffeas \storeregister[22][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][22] .is_wysiwyg = "true";
defparam \storeregister[22][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N26
cycloneive_lcell_comb \Mux9~3 (
// Equation(s):
// \Mux9~3_combout  = (\Mux9~2_combout  & (((\storeregister[30][22]~q )) # (!temp_imemload_output_23))) # (!\Mux9~2_combout  & (temp_imemload_output_23 & ((\storeregister[22][22]~q ))))

	.dataa(\Mux9~2_combout ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[30][22]~q ),
	.datad(\storeregister[22][22]~q ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~3 .lut_mask = 16'hE6A2;
defparam \Mux9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N15
dffeas \storeregister[28][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][22] .is_wysiwyg = "true";
defparam \storeregister[28][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y35_N5
dffeas \storeregister[16][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][22] .is_wysiwyg = "true";
defparam \storeregister[16][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N24
cycloneive_lcell_comb \storeregister[24][22]~feeder (
// Equation(s):
// \storeregister[24][22]~feeder_combout  = Mux9

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux9),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[24][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][22]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[24][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N25
dffeas \storeregister[24][22] (
	.clk(!CLK),
	.d(\storeregister[24][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][22] .is_wysiwyg = "true";
defparam \storeregister[24][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N4
cycloneive_lcell_comb \Mux9~4 (
// Equation(s):
// \Mux9~4_combout  = (temp_imemload_output_23 & (temp_imemload_output_24)) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & ((\storeregister[24][22]~q ))) # (!temp_imemload_output_24 & (\storeregister[16][22]~q ))))

	.dataa(temp_imemload_output_23),
	.datab(temp_imemload_output_24),
	.datac(\storeregister[16][22]~q ),
	.datad(\storeregister[24][22]~q ),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~4 .lut_mask = 16'hDC98;
defparam \Mux9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N14
cycloneive_lcell_comb \Mux9~5 (
// Equation(s):
// \Mux9~5_combout  = (temp_imemload_output_23 & ((\Mux9~4_combout  & ((\storeregister[28][22]~q ))) # (!\Mux9~4_combout  & (\storeregister[20][22]~q )))) # (!temp_imemload_output_23 & (((\Mux9~4_combout ))))

	.dataa(\storeregister[20][22]~q ),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[28][22]~q ),
	.datad(\Mux9~4_combout ),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~5 .lut_mask = 16'hF388;
defparam \Mux9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N28
cycloneive_lcell_comb \Mux9~6 (
// Equation(s):
// \Mux9~6_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\Mux9~3_combout )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & ((\Mux9~5_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\Mux9~3_combout ),
	.datad(\Mux9~5_combout ),
	.cin(gnd),
	.combout(\Mux9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~6 .lut_mask = 16'hB9A8;
defparam \Mux9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N19
dffeas \storeregister[10][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][22] .is_wysiwyg = "true";
defparam \storeregister[10][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N18
cycloneive_lcell_comb \Mux9~10 (
// Equation(s):
// \Mux9~10_combout  = (temp_imemload_output_22 & (((\storeregister[10][22]~q ) # (temp_imemload_output_21)))) # (!temp_imemload_output_22 & (\storeregister[8][22]~q  & ((!temp_imemload_output_21))))

	.dataa(\storeregister[8][22]~q ),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[10][22]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux9~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~10 .lut_mask = 16'hCCE2;
defparam \Mux9~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N9
dffeas \storeregister[9][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][22] .is_wysiwyg = "true";
defparam \storeregister[9][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N23
dffeas \storeregister[11][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][22] .is_wysiwyg = "true";
defparam \storeregister[11][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N8
cycloneive_lcell_comb \Mux9~11 (
// Equation(s):
// \Mux9~11_combout  = (\Mux9~10_combout  & (((\storeregister[11][22]~q )) # (!temp_imemload_output_21))) # (!\Mux9~10_combout  & (temp_imemload_output_21 & (\storeregister[9][22]~q )))

	.dataa(\Mux9~10_combout ),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[9][22]~q ),
	.datad(\storeregister[11][22]~q ),
	.cin(gnd),
	.combout(\Mux9~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~11 .lut_mask = 16'hEA62;
defparam \Mux9~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N0
cycloneive_lcell_comb \storeregister[14][22]~feeder (
// Equation(s):
// \storeregister[14][22]~feeder_combout  = Mux9

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux9),
	.cin(gnd),
	.combout(\storeregister[14][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][22]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[14][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N1
dffeas \storeregister[14][22] (
	.clk(!CLK),
	.d(\storeregister[14][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][22] .is_wysiwyg = "true";
defparam \storeregister[14][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N23
dffeas \storeregister[15][22] (
	.clk(!CLK),
	.d(Mux9),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][22] .is_wysiwyg = "true";
defparam \storeregister[15][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N17
dffeas \storeregister[13][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][22] .is_wysiwyg = "true";
defparam \storeregister[13][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N11
dffeas \storeregister[12][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][22] .is_wysiwyg = "true";
defparam \storeregister[12][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N16
cycloneive_lcell_comb \Mux9~17 (
// Equation(s):
// \Mux9~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][22]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[12][22]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[13][22]~q ),
	.datad(\storeregister[12][22]~q ),
	.cin(gnd),
	.combout(\Mux9~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~17 .lut_mask = 16'hB9A8;
defparam \Mux9~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N18
cycloneive_lcell_comb \Mux9~18 (
// Equation(s):
// \Mux9~18_combout  = (temp_imemload_output_22 & ((\Mux9~17_combout  & ((\storeregister[15][22]~q ))) # (!\Mux9~17_combout  & (\storeregister[14][22]~q )))) # (!temp_imemload_output_22 & (((\Mux9~17_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[14][22]~q ),
	.datac(\storeregister[15][22]~q ),
	.datad(\Mux9~17_combout ),
	.cin(gnd),
	.combout(\Mux9~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~18 .lut_mask = 16'hF588;
defparam \Mux9~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y41_N23
dffeas \storeregister[4][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][22] .is_wysiwyg = "true";
defparam \storeregister[4][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y41_N1
dffeas \storeregister[5][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][22] .is_wysiwyg = "true";
defparam \storeregister[5][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N22
cycloneive_lcell_comb \Mux9~12 (
// Equation(s):
// \Mux9~12_combout  = (temp_imemload_output_22 & (temp_imemload_output_21)) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & ((\storeregister[5][22]~q ))) # (!temp_imemload_output_21 & (\storeregister[4][22]~q ))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[4][22]~q ),
	.datad(\storeregister[5][22]~q ),
	.cin(gnd),
	.combout(\Mux9~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~12 .lut_mask = 16'hDC98;
defparam \Mux9~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N29
dffeas \storeregister[7][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][22] .is_wysiwyg = "true";
defparam \storeregister[7][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N3
dffeas \storeregister[6][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][22] .is_wysiwyg = "true";
defparam \storeregister[6][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N28
cycloneive_lcell_comb \Mux9~13 (
// Equation(s):
// \Mux9~13_combout  = (temp_imemload_output_22 & ((\Mux9~12_combout  & (\storeregister[7][22]~q )) # (!\Mux9~12_combout  & ((\storeregister[6][22]~q ))))) # (!temp_imemload_output_22 & (\Mux9~12_combout ))

	.dataa(temp_imemload_output_22),
	.datab(\Mux9~12_combout ),
	.datac(\storeregister[7][22]~q ),
	.datad(\storeregister[6][22]~q ),
	.cin(gnd),
	.combout(\Mux9~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~13 .lut_mask = 16'hE6C4;
defparam \Mux9~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N3
dffeas \storeregister[2][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][22] .is_wysiwyg = "true";
defparam \storeregister[2][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N16
cycloneive_lcell_comb \Mux9~15 (
// Equation(s):
// \Mux9~15_combout  = (\Mux9~14_combout ) # ((!temp_imemload_output_21 & (temp_imemload_output_22 & \storeregister[2][22]~q )))

	.dataa(\Mux9~14_combout ),
	.datab(temp_imemload_output_21),
	.datac(temp_imemload_output_22),
	.datad(\storeregister[2][22]~q ),
	.cin(gnd),
	.combout(\Mux9~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~15 .lut_mask = 16'hBAAA;
defparam \Mux9~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N14
cycloneive_lcell_comb \Mux9~16 (
// Equation(s):
// \Mux9~16_combout  = (temp_imemload_output_24 & (((temp_imemload_output_23)))) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\Mux9~13_combout )) # (!temp_imemload_output_23 & ((\Mux9~15_combout )))))

	.dataa(temp_imemload_output_24),
	.datab(\Mux9~13_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux9~15_combout ),
	.cin(gnd),
	.combout(\Mux9~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~16 .lut_mask = 16'hE5E0;
defparam \Mux9~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N16
cycloneive_lcell_comb \storeregister[24][21]~feeder (
// Equation(s):
// \storeregister[24][21]~feeder_combout  = Mux10

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux10),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[24][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][21]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[24][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N17
dffeas \storeregister[24][21] (
	.clk(!CLK),
	.d(\storeregister[24][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][21] .is_wysiwyg = "true";
defparam \storeregister[24][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N25
dffeas \storeregister[28][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][21] .is_wysiwyg = "true";
defparam \storeregister[28][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N24
cycloneive_lcell_comb \Mux10~5 (
// Equation(s):
// \Mux10~5_combout  = (\Mux10~4_combout  & (((\storeregister[28][21]~q ) # (!temp_imemload_output_24)))) # (!\Mux10~4_combout  & (\storeregister[24][21]~q  & ((temp_imemload_output_24))))

	.dataa(\Mux10~4_combout ),
	.datab(\storeregister[24][21]~q ),
	.datac(\storeregister[28][21]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~5 .lut_mask = 16'hE4AA;
defparam \Mux10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N1
dffeas \storeregister[22][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][21] .is_wysiwyg = "true";
defparam \storeregister[22][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N27
dffeas \storeregister[18][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][21] .is_wysiwyg = "true";
defparam \storeregister[18][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N0
cycloneive_lcell_comb \Mux10~2 (
// Equation(s):
// \Mux10~2_combout  = (temp_imemload_output_24 & (temp_imemload_output_23)) # (!temp_imemload_output_24 & ((temp_imemload_output_23 & (\storeregister[22][21]~q )) # (!temp_imemload_output_23 & ((\storeregister[18][21]~q )))))

	.dataa(temp_imemload_output_24),
	.datab(temp_imemload_output_23),
	.datac(\storeregister[22][21]~q ),
	.datad(\storeregister[18][21]~q ),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~2 .lut_mask = 16'hD9C8;
defparam \Mux10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N17
dffeas \storeregister[26][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][21] .is_wysiwyg = "true";
defparam \storeregister[26][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N16
cycloneive_lcell_comb \Mux10~3 (
// Equation(s):
// \Mux10~3_combout  = (\Mux10~2_combout  & ((\storeregister[30][21]~q ) # ((!temp_imemload_output_24)))) # (!\Mux10~2_combout  & (((\storeregister[26][21]~q  & temp_imemload_output_24))))

	.dataa(\storeregister[30][21]~q ),
	.datab(\Mux10~2_combout ),
	.datac(\storeregister[26][21]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~3 .lut_mask = 16'hB8CC;
defparam \Mux10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N12
cycloneive_lcell_comb \Mux10~6 (
// Equation(s):
// \Mux10~6_combout  = (temp_imemload_output_21 & (((temp_imemload_output_22)))) # (!temp_imemload_output_21 & ((temp_imemload_output_22 & ((\Mux10~3_combout ))) # (!temp_imemload_output_22 & (\Mux10~5_combout ))))

	.dataa(\Mux10~5_combout ),
	.datab(temp_imemload_output_21),
	.datac(\Mux10~3_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~6 .lut_mask = 16'hFC22;
defparam \Mux10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N23
dffeas \storeregister[21][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][21] .is_wysiwyg = "true";
defparam \storeregister[21][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N29
dffeas \storeregister[29][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[29][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[29][21] .is_wysiwyg = "true";
defparam \storeregister[29][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N24
cycloneive_lcell_comb \storeregister[25][21]~feeder (
// Equation(s):
// \storeregister[25][21]~feeder_combout  = Mux10

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux10),
	.cin(gnd),
	.combout(\storeregister[25][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[25][21]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[25][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N25
dffeas \storeregister[25][21] (
	.clk(!CLK),
	.d(\storeregister[25][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][21] .is_wysiwyg = "true";
defparam \storeregister[25][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N7
dffeas \storeregister[17][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][21] .is_wysiwyg = "true";
defparam \storeregister[17][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N6
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[25][21]~q )) # (!temp_imemload_output_24 & ((\storeregister[17][21]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[25][21]~q ),
	.datac(\storeregister[17][21]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hEE50;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N28
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (temp_imemload_output_23 & ((\Mux10~0_combout  & ((\storeregister[29][21]~q ))) # (!\Mux10~0_combout  & (\storeregister[21][21]~q )))) # (!temp_imemload_output_23 & (((\Mux10~0_combout ))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[21][21]~q ),
	.datac(\storeregister[29][21]~q ),
	.datad(\Mux10~0_combout ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hF588;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N18
cycloneive_lcell_comb \storeregister[27][21]~feeder (
// Equation(s):
// \storeregister[27][21]~feeder_combout  = Mux10

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux10),
	.cin(gnd),
	.combout(\storeregister[27][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][21]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[27][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N19
dffeas \storeregister[27][21] (
	.clk(!CLK),
	.d(\storeregister[27][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][21] .is_wysiwyg = "true";
defparam \storeregister[27][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N6
cycloneive_lcell_comb \storeregister[19][21]~feeder (
// Equation(s):
// \storeregister[19][21]~feeder_combout  = Mux10

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux10),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[19][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[19][21]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[19][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N7
dffeas \storeregister[19][21] (
	.clk(!CLK),
	.d(\storeregister[19][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][21] .is_wysiwyg = "true";
defparam \storeregister[19][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N8
cycloneive_lcell_comb \Mux10~7 (
// Equation(s):
// \Mux10~7_combout  = (temp_imemload_output_23 & (((temp_imemload_output_24)))) # (!temp_imemload_output_23 & ((temp_imemload_output_24 & (\storeregister[27][21]~q )) # (!temp_imemload_output_24 & ((\storeregister[19][21]~q )))))

	.dataa(temp_imemload_output_23),
	.datab(\storeregister[27][21]~q ),
	.datac(\storeregister[19][21]~q ),
	.datad(temp_imemload_output_24),
	.cin(gnd),
	.combout(\Mux10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~7 .lut_mask = 16'hEE50;
defparam \Mux10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N13
dffeas \storeregister[31][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[31][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[31][21] .is_wysiwyg = "true";
defparam \storeregister[31][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N1
dffeas \storeregister[23][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][21] .is_wysiwyg = "true";
defparam \storeregister[23][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N12
cycloneive_lcell_comb \Mux10~8 (
// Equation(s):
// \Mux10~8_combout  = (temp_imemload_output_23 & ((\Mux10~7_combout  & (\storeregister[31][21]~q )) # (!\Mux10~7_combout  & ((\storeregister[23][21]~q ))))) # (!temp_imemload_output_23 & (\Mux10~7_combout ))

	.dataa(temp_imemload_output_23),
	.datab(\Mux10~7_combout ),
	.datac(\storeregister[31][21]~q ),
	.datad(\storeregister[23][21]~q ),
	.cin(gnd),
	.combout(\Mux10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~8 .lut_mask = 16'hE6C4;
defparam \Mux10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N31
dffeas \storeregister[8][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][21] .is_wysiwyg = "true";
defparam \storeregister[8][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N1
dffeas \storeregister[10][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][21] .is_wysiwyg = "true";
defparam \storeregister[10][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N30
cycloneive_lcell_comb \Mux10~12 (
// Equation(s):
// \Mux10~12_combout  = (temp_imemload_output_22 & ((temp_imemload_output_21) # ((\storeregister[10][21]~q )))) # (!temp_imemload_output_22 & (!temp_imemload_output_21 & (\storeregister[8][21]~q )))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[8][21]~q ),
	.datad(\storeregister[10][21]~q ),
	.cin(gnd),
	.combout(\Mux10~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~12 .lut_mask = 16'hBA98;
defparam \Mux10~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N27
dffeas \storeregister[11][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][21] .is_wysiwyg = "true";
defparam \storeregister[11][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N26
cycloneive_lcell_comb \Mux10~13 (
// Equation(s):
// \Mux10~13_combout  = (\Mux10~12_combout  & (((\storeregister[11][21]~q ) # (!temp_imemload_output_21)))) # (!\Mux10~12_combout  & (\storeregister[9][21]~q  & ((temp_imemload_output_21))))

	.dataa(\storeregister[9][21]~q ),
	.datab(\Mux10~12_combout ),
	.datac(\storeregister[11][21]~q ),
	.datad(temp_imemload_output_21),
	.cin(gnd),
	.combout(\Mux10~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~13 .lut_mask = 16'hE2CC;
defparam \Mux10~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N1
dffeas \storeregister[3][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][21] .is_wysiwyg = "true";
defparam \storeregister[3][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N3
dffeas \storeregister[1][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][21] .is_wysiwyg = "true";
defparam \storeregister[1][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N0
cycloneive_lcell_comb \Mux10~14 (
// Equation(s):
// \Mux10~14_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22 & (\storeregister[3][21]~q )) # (!temp_imemload_output_22 & ((\storeregister[1][21]~q )))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[3][21]~q ),
	.datad(\storeregister[1][21]~q ),
	.cin(gnd),
	.combout(\Mux10~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~14 .lut_mask = 16'hA280;
defparam \Mux10~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N20
cycloneive_lcell_comb \Mux10~15 (
// Equation(s):
// \Mux10~15_combout  = (\Mux10~14_combout ) # ((\storeregister[2][21]~q  & (!temp_imemload_output_21 & temp_imemload_output_22)))

	.dataa(\storeregister[2][21]~q ),
	.datab(temp_imemload_output_21),
	.datac(\Mux10~14_combout ),
	.datad(temp_imemload_output_22),
	.cin(gnd),
	.combout(\Mux10~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~15 .lut_mask = 16'hF2F0;
defparam \Mux10~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N10
cycloneive_lcell_comb \Mux10~16 (
// Equation(s):
// \Mux10~16_combout  = (temp_imemload_output_24 & ((\Mux10~13_combout ) # ((temp_imemload_output_23)))) # (!temp_imemload_output_24 & (((!temp_imemload_output_23 & \Mux10~15_combout ))))

	.dataa(temp_imemload_output_24),
	.datab(\Mux10~13_combout ),
	.datac(temp_imemload_output_23),
	.datad(\Mux10~15_combout ),
	.cin(gnd),
	.combout(\Mux10~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~16 .lut_mask = 16'hADA8;
defparam \Mux10~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N26
cycloneive_lcell_comb \storeregister[15][21]~feeder (
// Equation(s):
// \storeregister[15][21]~feeder_combout  = Mux10

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux10),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[15][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[15][21]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[15][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N27
dffeas \storeregister[15][21] (
	.clk(!CLK),
	.d(\storeregister[15][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[15][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[15][21] .is_wysiwyg = "true";
defparam \storeregister[15][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N1
dffeas \storeregister[13][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][21] .is_wysiwyg = "true";
defparam \storeregister[13][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N19
dffeas \storeregister[12][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][21] .is_wysiwyg = "true";
defparam \storeregister[12][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N0
cycloneive_lcell_comb \Mux10~17 (
// Equation(s):
// \Mux10~17_combout  = (temp_imemload_output_21 & ((temp_imemload_output_22) # ((\storeregister[13][21]~q )))) # (!temp_imemload_output_21 & (!temp_imemload_output_22 & ((\storeregister[12][21]~q ))))

	.dataa(temp_imemload_output_21),
	.datab(temp_imemload_output_22),
	.datac(\storeregister[13][21]~q ),
	.datad(\storeregister[12][21]~q ),
	.cin(gnd),
	.combout(\Mux10~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~17 .lut_mask = 16'hB9A8;
defparam \Mux10~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N16
cycloneive_lcell_comb \storeregister[14][21]~feeder (
// Equation(s):
// \storeregister[14][21]~feeder_combout  = Mux10

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux10),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[14][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[14][21]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[14][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N17
dffeas \storeregister[14][21] (
	.clk(!CLK),
	.d(\storeregister[14][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[14][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[14][21] .is_wysiwyg = "true";
defparam \storeregister[14][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N24
cycloneive_lcell_comb \Mux10~18 (
// Equation(s):
// \Mux10~18_combout  = (temp_imemload_output_22 & ((\Mux10~17_combout  & (\storeregister[15][21]~q )) # (!\Mux10~17_combout  & ((\storeregister[14][21]~q ))))) # (!temp_imemload_output_22 & (((\Mux10~17_combout ))))

	.dataa(\storeregister[15][21]~q ),
	.datab(temp_imemload_output_22),
	.datac(\Mux10~17_combout ),
	.datad(\storeregister[14][21]~q ),
	.cin(gnd),
	.combout(\Mux10~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~18 .lut_mask = 16'hBCB0;
defparam \Mux10~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N5
dffeas \storeregister[7][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[7][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[7][21] .is_wysiwyg = "true";
defparam \storeregister[7][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N23
dffeas \storeregister[6][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][21] .is_wysiwyg = "true";
defparam \storeregister[6][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y41_N25
dffeas \storeregister[5][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][21] .is_wysiwyg = "true";
defparam \storeregister[5][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y41_N7
dffeas \storeregister[4][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][21] .is_wysiwyg = "true";
defparam \storeregister[4][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N24
cycloneive_lcell_comb \Mux10~10 (
// Equation(s):
// \Mux10~10_combout  = (temp_imemload_output_22 & (temp_imemload_output_21)) # (!temp_imemload_output_22 & ((temp_imemload_output_21 & (\storeregister[5][21]~q )) # (!temp_imemload_output_21 & ((\storeregister[4][21]~q )))))

	.dataa(temp_imemload_output_22),
	.datab(temp_imemload_output_21),
	.datac(\storeregister[5][21]~q ),
	.datad(\storeregister[4][21]~q ),
	.cin(gnd),
	.combout(\Mux10~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~10 .lut_mask = 16'hD9C8;
defparam \Mux10~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N22
cycloneive_lcell_comb \Mux10~11 (
// Equation(s):
// \Mux10~11_combout  = (temp_imemload_output_22 & ((\Mux10~10_combout  & (\storeregister[7][21]~q )) # (!\Mux10~10_combout  & ((\storeregister[6][21]~q ))))) # (!temp_imemload_output_22 & (((\Mux10~10_combout ))))

	.dataa(temp_imemload_output_22),
	.datab(\storeregister[7][21]~q ),
	.datac(\storeregister[6][21]~q ),
	.datad(\Mux10~10_combout ),
	.cin(gnd),
	.combout(\Mux10~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~11 .lut_mask = 16'hDDA0;
defparam \Mux10~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N9
dffeas \storeregister[20][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][15] .is_wysiwyg = "true";
defparam \storeregister[20][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N11
dffeas \storeregister[16][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][15] .is_wysiwyg = "true";
defparam \storeregister[16][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N10
cycloneive_lcell_comb \Mux48~4 (
// Equation(s):
// \Mux48~4_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\storeregister[24][15]~q )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & (\storeregister[16][15]~q )))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[16][15]~q ),
	.datad(\storeregister[24][15]~q ),
	.cin(gnd),
	.combout(\Mux48~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~4 .lut_mask = 16'hBA98;
defparam \Mux48~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N0
cycloneive_lcell_comb \Mux48~5 (
// Equation(s):
// \Mux48~5_combout  = (temp_imemload_output_18 & ((\Mux48~4_combout  & ((\storeregister[28][15]~q ))) # (!\Mux48~4_combout  & (\storeregister[20][15]~q )))) # (!temp_imemload_output_18 & (((\Mux48~4_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[20][15]~q ),
	.datac(\storeregister[28][15]~q ),
	.datad(\Mux48~4_combout ),
	.cin(gnd),
	.combout(\Mux48~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~5 .lut_mask = 16'hF588;
defparam \Mux48~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N6
cycloneive_lcell_comb \Mux48~3 (
// Equation(s):
// \Mux48~3_combout  = (\Mux48~2_combout  & (((\storeregister[30][15]~q ) # (!temp_imemload_output_18)))) # (!\Mux48~2_combout  & (\storeregister[22][15]~q  & ((temp_imemload_output_18))))

	.dataa(\Mux48~2_combout ),
	.datab(\storeregister[22][15]~q ),
	.datac(\storeregister[30][15]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux48~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~3 .lut_mask = 16'hE4AA;
defparam \Mux48~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N12
cycloneive_lcell_comb \Mux48~6 (
// Equation(s):
// \Mux48~6_combout  = (temp_imemload_output_17 & ((temp_imemload_output_16) # ((\Mux48~3_combout )))) # (!temp_imemload_output_17 & (!temp_imemload_output_16 & (\Mux48~5_combout )))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\Mux48~5_combout ),
	.datad(\Mux48~3_combout ),
	.cin(gnd),
	.combout(\Mux48~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~6 .lut_mask = 16'hBA98;
defparam \Mux48~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N6
cycloneive_lcell_comb \storeregister[19][15]~feeder (
// Equation(s):
// \storeregister[19][15]~feeder_combout  = Mux16

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux16),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[19][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[19][15]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[19][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N7
dffeas \storeregister[19][15] (
	.clk(!CLK),
	.d(\storeregister[19][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][15] .is_wysiwyg = "true";
defparam \storeregister[19][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N14
cycloneive_lcell_comb \Mux48~7 (
// Equation(s):
// \Mux48~7_combout  = (temp_imemload_output_18 & ((\storeregister[23][15]~q ) # ((temp_imemload_output_19)))) # (!temp_imemload_output_18 & (((\storeregister[19][15]~q  & !temp_imemload_output_19))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[23][15]~q ),
	.datac(\storeregister[19][15]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux48~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~7 .lut_mask = 16'hAAD8;
defparam \Mux48~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N0
cycloneive_lcell_comb \Mux48~8 (
// Equation(s):
// \Mux48~8_combout  = (temp_imemload_output_19 & ((\Mux48~7_combout  & ((\storeregister[31][15]~q ))) # (!\Mux48~7_combout  & (\storeregister[27][15]~q )))) # (!temp_imemload_output_19 & (\Mux48~7_combout ))

	.dataa(temp_imemload_output_19),
	.datab(\Mux48~7_combout ),
	.datac(\storeregister[27][15]~q ),
	.datad(\storeregister[31][15]~q ),
	.cin(gnd),
	.combout(\Mux48~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~8 .lut_mask = 16'hEC64;
defparam \Mux48~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N24
cycloneive_lcell_comb \Mux48~0 (
// Equation(s):
// \Mux48~0_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[21][15]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[17][15]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[21][15]~q ),
	.datad(\storeregister[17][15]~q ),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~0 .lut_mask = 16'hB9A8;
defparam \Mux48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N22
cycloneive_lcell_comb \Mux48~1 (
// Equation(s):
// \Mux48~1_combout  = (\Mux48~0_combout  & ((\storeregister[29][15]~q ) # ((!temp_imemload_output_19)))) # (!\Mux48~0_combout  & (((temp_imemload_output_19 & \storeregister[25][15]~q ))))

	.dataa(\Mux48~0_combout ),
	.datab(\storeregister[29][15]~q ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[25][15]~q ),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~1 .lut_mask = 16'hDA8A;
defparam \Mux48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N26
cycloneive_lcell_comb \Mux48~17 (
// Equation(s):
// \Mux48~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][15]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][15]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[12][15]~q ),
	.datad(\storeregister[13][15]~q ),
	.cin(gnd),
	.combout(\Mux48~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~17 .lut_mask = 16'hDC98;
defparam \Mux48~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N12
cycloneive_lcell_comb \Mux48~18 (
// Equation(s):
// \Mux48~18_combout  = (\Mux48~17_combout  & ((\storeregister[15][15]~q ) # ((!temp_imemload_output_17)))) # (!\Mux48~17_combout  & (((temp_imemload_output_17 & \storeregister[14][15]~q ))))

	.dataa(\Mux48~17_combout ),
	.datab(\storeregister[15][15]~q ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[14][15]~q ),
	.cin(gnd),
	.combout(\Mux48~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~18 .lut_mask = 16'hDA8A;
defparam \Mux48~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N2
cycloneive_lcell_comb \Mux48~12 (
// Equation(s):
// \Mux48~12_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[5][15]~q )) # (!temp_imemload_output_16 & ((\storeregister[4][15]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[5][15]~q ),
	.datac(\storeregister[4][15]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux48~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~12 .lut_mask = 16'hEE50;
defparam \Mux48~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N22
cycloneive_lcell_comb \Mux48~13 (
// Equation(s):
// \Mux48~13_combout  = (temp_imemload_output_17 & ((\Mux48~12_combout  & ((\storeregister[7][15]~q ))) # (!\Mux48~12_combout  & (\storeregister[6][15]~q )))) # (!temp_imemload_output_17 & (((\Mux48~12_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[6][15]~q ),
	.datac(\storeregister[7][15]~q ),
	.datad(\Mux48~12_combout ),
	.cin(gnd),
	.combout(\Mux48~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~13 .lut_mask = 16'hF588;
defparam \Mux48~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N8
cycloneive_lcell_comb \Mux48~14 (
// Equation(s):
// \Mux48~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][15]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][15]~q )))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[3][15]~q ),
	.datad(\storeregister[1][15]~q ),
	.cin(gnd),
	.combout(\Mux48~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~14 .lut_mask = 16'hA280;
defparam \Mux48~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N20
cycloneive_lcell_comb \Mux48~15 (
// Equation(s):
// \Mux48~15_combout  = (\Mux48~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][15]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux48~14_combout ),
	.datac(\storeregister[2][15]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux48~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~15 .lut_mask = 16'hCCEC;
defparam \Mux48~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N26
cycloneive_lcell_comb \Mux48~16 (
// Equation(s):
// \Mux48~16_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\Mux48~13_combout )) # (!temp_imemload_output_18 & ((\Mux48~15_combout )))))

	.dataa(\Mux48~13_combout ),
	.datab(\Mux48~15_combout ),
	.datac(temp_imemload_output_19),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux48~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~16 .lut_mask = 16'hFA0C;
defparam \Mux48~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N31
dffeas \storeregister[10][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][15] .is_wysiwyg = "true";
defparam \storeregister[10][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N17
dffeas \storeregister[8][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][15] .is_wysiwyg = "true";
defparam \storeregister[8][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N30
cycloneive_lcell_comb \Mux48~10 (
// Equation(s):
// \Mux48~10_combout  = (temp_imemload_output_17 & ((temp_imemload_output_16) # ((\storeregister[10][15]~q )))) # (!temp_imemload_output_17 & (!temp_imemload_output_16 & ((\storeregister[8][15]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[10][15]~q ),
	.datad(\storeregister[8][15]~q ),
	.cin(gnd),
	.combout(\Mux48~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~10 .lut_mask = 16'hB9A8;
defparam \Mux48~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N0
cycloneive_lcell_comb \Mux48~11 (
// Equation(s):
// \Mux48~11_combout  = (\Mux48~10_combout  & ((\storeregister[11][15]~q ) # ((!temp_imemload_output_16)))) # (!\Mux48~10_combout  & (((\storeregister[9][15]~q  & temp_imemload_output_16))))

	.dataa(\storeregister[11][15]~q ),
	.datab(\Mux48~10_combout ),
	.datac(\storeregister[9][15]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux48~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~11 .lut_mask = 16'hB8CC;
defparam \Mux48~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N14
cycloneive_lcell_comb \Mux51~7 (
// Equation(s):
// \Mux51~7_combout  = (temp_imemload_output_19 & ((\storeregister[27][12]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((!temp_imemload_output_18 & \storeregister[19][12]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[27][12]~q ),
	.datac(temp_imemload_output_18),
	.datad(\storeregister[19][12]~q ),
	.cin(gnd),
	.combout(\Mux51~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~7 .lut_mask = 16'hADA8;
defparam \Mux51~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N14
cycloneive_lcell_comb \Mux51~8 (
// Equation(s):
// \Mux51~8_combout  = (\Mux51~7_combout  & (((\storeregister[31][12]~q )) # (!temp_imemload_output_18))) # (!\Mux51~7_combout  & (temp_imemload_output_18 & (\storeregister[23][12]~q )))

	.dataa(\Mux51~7_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[23][12]~q ),
	.datad(\storeregister[31][12]~q ),
	.cin(gnd),
	.combout(\Mux51~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~8 .lut_mask = 16'hEA62;
defparam \Mux51~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N10
cycloneive_lcell_comb \Mux51~0 (
// Equation(s):
// \Mux51~0_combout  = (temp_imemload_output_19 & ((\storeregister[25][12]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\storeregister[17][12]~q  & !temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[25][12]~q ),
	.datac(\storeregister[17][12]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~0 .lut_mask = 16'hAAD8;
defparam \Mux51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N0
cycloneive_lcell_comb \Mux51~1 (
// Equation(s):
// \Mux51~1_combout  = (temp_imemload_output_18 & ((\Mux51~0_combout  & ((\storeregister[29][12]~q ))) # (!\Mux51~0_combout  & (\storeregister[21][12]~q )))) # (!temp_imemload_output_18 & (\Mux51~0_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux51~0_combout ),
	.datac(\storeregister[21][12]~q ),
	.datad(\storeregister[29][12]~q ),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~1 .lut_mask = 16'hEC64;
defparam \Mux51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N4
cycloneive_lcell_comb \Mux51~2 (
// Equation(s):
// \Mux51~2_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[22][12]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[18][12]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[18][12]~q ),
	.datad(\storeregister[22][12]~q ),
	.cin(gnd),
	.combout(\Mux51~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~2 .lut_mask = 16'hBA98;
defparam \Mux51~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N10
cycloneive_lcell_comb \Mux51~3 (
// Equation(s):
// \Mux51~3_combout  = (\Mux51~2_combout  & ((\storeregister[30][12]~q ) # ((!temp_imemload_output_19)))) # (!\Mux51~2_combout  & (((\storeregister[26][12]~q  & temp_imemload_output_19))))

	.dataa(\storeregister[30][12]~q ),
	.datab(\Mux51~2_combout ),
	.datac(\storeregister[26][12]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux51~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~3 .lut_mask = 16'hB8CC;
defparam \Mux51~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N28
cycloneive_lcell_comb \Mux51~4 (
// Equation(s):
// \Mux51~4_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[20][12]~q ))) # (!temp_imemload_output_18 & (\storeregister[16][12]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[16][12]~q ),
	.datac(\storeregister[20][12]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux51~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~4 .lut_mask = 16'hFA44;
defparam \Mux51~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N0
cycloneive_lcell_comb \Mux51~5 (
// Equation(s):
// \Mux51~5_combout  = (temp_imemload_output_19 & ((\Mux51~4_combout  & ((\storeregister[28][12]~q ))) # (!\Mux51~4_combout  & (\storeregister[24][12]~q )))) # (!temp_imemload_output_19 & (((\Mux51~4_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[24][12]~q ),
	.datac(\Mux51~4_combout ),
	.datad(\storeregister[28][12]~q ),
	.cin(gnd),
	.combout(\Mux51~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~5 .lut_mask = 16'hF858;
defparam \Mux51~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N8
cycloneive_lcell_comb \Mux51~6 (
// Equation(s):
// \Mux51~6_combout  = (temp_imemload_output_17 & ((\Mux51~3_combout ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((\Mux51~5_combout  & !temp_imemload_output_16))))

	.dataa(\Mux51~3_combout ),
	.datab(\Mux51~5_combout ),
	.datac(temp_imemload_output_17),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux51~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~6 .lut_mask = 16'hF0AC;
defparam \Mux51~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N24
cycloneive_lcell_comb \Mux51~12 (
// Equation(s):
// \Mux51~12_combout  = (temp_imemload_output_17 & ((temp_imemload_output_16) # ((\storeregister[10][12]~q )))) # (!temp_imemload_output_17 & (!temp_imemload_output_16 & (\storeregister[8][12]~q )))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[8][12]~q ),
	.datad(\storeregister[10][12]~q ),
	.cin(gnd),
	.combout(\Mux51~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~12 .lut_mask = 16'hBA98;
defparam \Mux51~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N20
cycloneive_lcell_comb \Mux51~13 (
// Equation(s):
// \Mux51~13_combout  = (temp_imemload_output_16 & ((\Mux51~12_combout  & ((\storeregister[11][12]~q ))) # (!\Mux51~12_combout  & (\storeregister[9][12]~q )))) # (!temp_imemload_output_16 & (((\Mux51~12_combout ))))

	.dataa(\storeregister[9][12]~q ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[11][12]~q ),
	.datad(\Mux51~12_combout ),
	.cin(gnd),
	.combout(\Mux51~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~13 .lut_mask = 16'hF388;
defparam \Mux51~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N2
cycloneive_lcell_comb \Mux51~14 (
// Equation(s):
// \Mux51~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[3][12]~q ))) # (!temp_imemload_output_17 & (\storeregister[1][12]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[1][12]~q ),
	.datad(\storeregister[3][12]~q ),
	.cin(gnd),
	.combout(\Mux51~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~14 .lut_mask = 16'hA820;
defparam \Mux51~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N18
cycloneive_lcell_comb \Mux51~15 (
// Equation(s):
// \Mux51~15_combout  = (\Mux51~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][12]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[2][12]~q ),
	.datac(\Mux51~14_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux51~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~15 .lut_mask = 16'hF0F8;
defparam \Mux51~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N8
cycloneive_lcell_comb \Mux51~16 (
// Equation(s):
// \Mux51~16_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\Mux51~13_combout )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & ((\Mux51~15_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\Mux51~13_combout ),
	.datad(\Mux51~15_combout ),
	.cin(gnd),
	.combout(\Mux51~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~16 .lut_mask = 16'hB9A8;
defparam \Mux51~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N28
cycloneive_lcell_comb \Mux51~17 (
// Equation(s):
// \Mux51~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[13][12]~q )) # (!temp_imemload_output_16 & ((\storeregister[12][12]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[13][12]~q ),
	.datad(\storeregister[12][12]~q ),
	.cin(gnd),
	.combout(\Mux51~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~17 .lut_mask = 16'hD9C8;
defparam \Mux51~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N22
cycloneive_lcell_comb \Mux51~18 (
// Equation(s):
// \Mux51~18_combout  = (\Mux51~17_combout  & (((\storeregister[15][12]~q )) # (!temp_imemload_output_17))) # (!\Mux51~17_combout  & (temp_imemload_output_17 & ((\storeregister[14][12]~q ))))

	.dataa(\Mux51~17_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[15][12]~q ),
	.datad(\storeregister[14][12]~q ),
	.cin(gnd),
	.combout(\Mux51~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~18 .lut_mask = 16'hE6A2;
defparam \Mux51~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y42_N19
dffeas \storeregister[4][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][12] .is_wysiwyg = "true";
defparam \storeregister[4][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y42_N21
dffeas \storeregister[5][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][12] .is_wysiwyg = "true";
defparam \storeregister[5][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N20
cycloneive_lcell_comb \Mux51~10 (
// Equation(s):
// \Mux51~10_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[5][12]~q ))) # (!temp_imemload_output_16 & (\storeregister[4][12]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[4][12]~q ),
	.datac(\storeregister[5][12]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux51~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~10 .lut_mask = 16'hFA44;
defparam \Mux51~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N20
cycloneive_lcell_comb \Mux51~11 (
// Equation(s):
// \Mux51~11_combout  = (temp_imemload_output_17 & ((\Mux51~10_combout  & (\storeregister[7][12]~q )) # (!\Mux51~10_combout  & ((\storeregister[6][12]~q ))))) # (!temp_imemload_output_17 & (((\Mux51~10_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[7][12]~q ),
	.datac(\storeregister[6][12]~q ),
	.datad(\Mux51~10_combout ),
	.cin(gnd),
	.combout(\Mux51~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~11 .lut_mask = 16'hDDA0;
defparam \Mux51~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N13
dffeas \storeregister[22][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][27] .is_wysiwyg = "true";
defparam \storeregister[22][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N27
dffeas \storeregister[18][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][27] .is_wysiwyg = "true";
defparam \storeregister[18][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N26
cycloneive_lcell_comb \Mux36~2 (
// Equation(s):
// \Mux36~2_combout  = (temp_imemload_output_18 & ((\storeregister[22][27]~q ) # ((temp_imemload_output_19)))) # (!temp_imemload_output_18 & (((\storeregister[18][27]~q  & !temp_imemload_output_19))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[22][27]~q ),
	.datac(\storeregister[18][27]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux36~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~2 .lut_mask = 16'hAAD8;
defparam \Mux36~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N0
cycloneive_lcell_comb \Mux36~3 (
// Equation(s):
// \Mux36~3_combout  = (temp_imemload_output_19 & ((\Mux36~2_combout  & (\storeregister[30][27]~q )) # (!\Mux36~2_combout  & ((\storeregister[26][27]~q ))))) # (!temp_imemload_output_19 & (((\Mux36~2_combout ))))

	.dataa(\storeregister[30][27]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[26][27]~q ),
	.datad(\Mux36~2_combout ),
	.cin(gnd),
	.combout(\Mux36~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~3 .lut_mask = 16'hBBC0;
defparam \Mux36~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N5
dffeas \storeregister[24][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][27] .is_wysiwyg = "true";
defparam \storeregister[24][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N6
cycloneive_lcell_comb \Mux36~4 (
// Equation(s):
// \Mux36~4_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[20][27]~q ))) # (!temp_imemload_output_18 & (\storeregister[16][27]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[16][27]~q ),
	.datad(\storeregister[20][27]~q ),
	.cin(gnd),
	.combout(\Mux36~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~4 .lut_mask = 16'hDC98;
defparam \Mux36~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N4
cycloneive_lcell_comb \Mux36~5 (
// Equation(s):
// \Mux36~5_combout  = (temp_imemload_output_19 & ((\Mux36~4_combout  & (\storeregister[28][27]~q )) # (!\Mux36~4_combout  & ((\storeregister[24][27]~q ))))) # (!temp_imemload_output_19 & (((\Mux36~4_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[28][27]~q ),
	.datac(\storeregister[24][27]~q ),
	.datad(\Mux36~4_combout ),
	.cin(gnd),
	.combout(\Mux36~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~5 .lut_mask = 16'hDDA0;
defparam \Mux36~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N2
cycloneive_lcell_comb \Mux36~6 (
// Equation(s):
// \Mux36~6_combout  = (temp_imemload_output_16 & (temp_imemload_output_17)) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\Mux36~3_combout )) # (!temp_imemload_output_17 & ((\Mux36~5_combout )))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\Mux36~3_combout ),
	.datad(\Mux36~5_combout ),
	.cin(gnd),
	.combout(\Mux36~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~6 .lut_mask = 16'hD9C8;
defparam \Mux36~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N28
cycloneive_lcell_comb \Mux36~0 (
// Equation(s):
// \Mux36~0_combout  = (temp_imemload_output_19 & (((\storeregister[25][27]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[17][27]~q  & ((!temp_imemload_output_18))))

	.dataa(\storeregister[17][27]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[25][27]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~0 .lut_mask = 16'hCCE2;
defparam \Mux36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N18
cycloneive_lcell_comb \Mux36~1 (
// Equation(s):
// \Mux36~1_combout  = (temp_imemload_output_18 & ((\Mux36~0_combout  & ((\storeregister[29][27]~q ))) # (!\Mux36~0_combout  & (\storeregister[21][27]~q )))) # (!temp_imemload_output_18 & (((\Mux36~0_combout ))))

	.dataa(\storeregister[21][27]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[29][27]~q ),
	.datad(\Mux36~0_combout ),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~1 .lut_mask = 16'hF388;
defparam \Mux36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N0
cycloneive_lcell_comb \Mux36~7 (
// Equation(s):
// \Mux36~7_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\storeregister[27][27]~q )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & ((\storeregister[19][27]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[27][27]~q ),
	.datad(\storeregister[19][27]~q ),
	.cin(gnd),
	.combout(\Mux36~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~7 .lut_mask = 16'hB9A8;
defparam \Mux36~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N22
cycloneive_lcell_comb \Mux36~8 (
// Equation(s):
// \Mux36~8_combout  = (\Mux36~7_combout  & (((\storeregister[31][27]~q )) # (!temp_imemload_output_18))) # (!\Mux36~7_combout  & (temp_imemload_output_18 & ((\storeregister[23][27]~q ))))

	.dataa(\Mux36~7_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[31][27]~q ),
	.datad(\storeregister[23][27]~q ),
	.cin(gnd),
	.combout(\Mux36~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~8 .lut_mask = 16'hE6A2;
defparam \Mux36~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N17
dffeas \storeregister[13][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][27] .is_wysiwyg = "true";
defparam \storeregister[13][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N16
cycloneive_lcell_comb \Mux36~17 (
// Equation(s):
// \Mux36~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[13][27]~q )) # (!temp_imemload_output_16 & ((\storeregister[12][27]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[13][27]~q ),
	.datad(\storeregister[12][27]~q ),
	.cin(gnd),
	.combout(\Mux36~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~17 .lut_mask = 16'hD9C8;
defparam \Mux36~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N4
cycloneive_lcell_comb \Mux36~18 (
// Equation(s):
// \Mux36~18_combout  = (\Mux36~17_combout  & (((\storeregister[15][27]~q )) # (!temp_imemload_output_17))) # (!\Mux36~17_combout  & (temp_imemload_output_17 & ((\storeregister[14][27]~q ))))

	.dataa(\Mux36~17_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[15][27]~q ),
	.datad(\storeregister[14][27]~q ),
	.cin(gnd),
	.combout(\Mux36~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~18 .lut_mask = 16'hE6A2;
defparam \Mux36~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N14
cycloneive_lcell_comb \Mux36~10 (
// Equation(s):
// \Mux36~10_combout  = (temp_imemload_output_16 & ((\storeregister[5][27]~q ) # ((temp_imemload_output_17)))) # (!temp_imemload_output_16 & (((\storeregister[4][27]~q  & !temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[5][27]~q ),
	.datac(\storeregister[4][27]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux36~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~10 .lut_mask = 16'hAAD8;
defparam \Mux36~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N4
cycloneive_lcell_comb \Mux36~11 (
// Equation(s):
// \Mux36~11_combout  = (\Mux36~10_combout  & (((\storeregister[7][27]~q )) # (!temp_imemload_output_17))) # (!\Mux36~10_combout  & (temp_imemload_output_17 & (\storeregister[6][27]~q )))

	.dataa(\Mux36~10_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[6][27]~q ),
	.datad(\storeregister[7][27]~q ),
	.cin(gnd),
	.combout(\Mux36~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~11 .lut_mask = 16'hEA62;
defparam \Mux36~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N10
cycloneive_lcell_comb \Mux36~15 (
// Equation(s):
// \Mux36~15_combout  = (\Mux36~14_combout ) # ((!temp_imemload_output_16 & (temp_imemload_output_17 & \storeregister[2][27]~q )))

	.dataa(\Mux36~14_combout ),
	.datab(temp_imemload_output_16),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[2][27]~q ),
	.cin(gnd),
	.combout(\Mux36~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~15 .lut_mask = 16'hBAAA;
defparam \Mux36~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N28
cycloneive_lcell_comb \Mux36~12 (
// Equation(s):
// \Mux36~12_combout  = (temp_imemload_output_17 & ((\storeregister[10][27]~q ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((\storeregister[8][27]~q  & !temp_imemload_output_16))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[10][27]~q ),
	.datac(\storeregister[8][27]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux36~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~12 .lut_mask = 16'hAAD8;
defparam \Mux36~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N14
cycloneive_lcell_comb \storeregister[9][27]~feeder (
// Equation(s):
// \storeregister[9][27]~feeder_combout  = Mux4

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux4),
	.cin(gnd),
	.combout(\storeregister[9][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[9][27]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[9][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N15
dffeas \storeregister[9][27] (
	.clk(!CLK),
	.d(\storeregister[9][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][27] .is_wysiwyg = "true";
defparam \storeregister[9][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N30
cycloneive_lcell_comb \Mux36~13 (
// Equation(s):
// \Mux36~13_combout  = (temp_imemload_output_16 & ((\Mux36~12_combout  & ((\storeregister[11][27]~q ))) # (!\Mux36~12_combout  & (\storeregister[9][27]~q )))) # (!temp_imemload_output_16 & (\Mux36~12_combout ))

	.dataa(temp_imemload_output_16),
	.datab(\Mux36~12_combout ),
	.datac(\storeregister[9][27]~q ),
	.datad(\storeregister[11][27]~q ),
	.cin(gnd),
	.combout(\Mux36~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~13 .lut_mask = 16'hEC64;
defparam \Mux36~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N20
cycloneive_lcell_comb \Mux36~16 (
// Equation(s):
// \Mux36~16_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18) # (\Mux36~13_combout )))) # (!temp_imemload_output_19 & (\Mux36~15_combout  & (!temp_imemload_output_18)))

	.dataa(\Mux36~15_combout ),
	.datab(temp_imemload_output_19),
	.datac(temp_imemload_output_18),
	.datad(\Mux36~13_combout ),
	.cin(gnd),
	.combout(\Mux36~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~16 .lut_mask = 16'hCEC2;
defparam \Mux36~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N30
cycloneive_lcell_comb \Mux45~7 (
// Equation(s):
// \Mux45~7_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[27][18]~q ))) # (!temp_imemload_output_19 & (\storeregister[19][18]~q ))))

	.dataa(\storeregister[19][18]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[27][18]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux45~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~7 .lut_mask = 16'hFC22;
defparam \Mux45~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N16
cycloneive_lcell_comb \Mux45~8 (
// Equation(s):
// \Mux45~8_combout  = (\Mux45~7_combout  & (((\storeregister[31][18]~q )) # (!temp_imemload_output_18))) # (!\Mux45~7_combout  & (temp_imemload_output_18 & (\storeregister[23][18]~q )))

	.dataa(\Mux45~7_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[23][18]~q ),
	.datad(\storeregister[31][18]~q ),
	.cin(gnd),
	.combout(\Mux45~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~8 .lut_mask = 16'hEA62;
defparam \Mux45~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N10
cycloneive_lcell_comb \Mux45~0 (
// Equation(s):
// \Mux45~0_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[25][18]~q ))) # (!temp_imemload_output_19 & (\storeregister[17][18]~q ))))

	.dataa(\storeregister[17][18]~q ),
	.datab(temp_imemload_output_18),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[25][18]~q ),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~0 .lut_mask = 16'hF2C2;
defparam \Mux45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N22
cycloneive_lcell_comb \Mux45~1 (
// Equation(s):
// \Mux45~1_combout  = (temp_imemload_output_18 & ((\Mux45~0_combout  & ((\storeregister[29][18]~q ))) # (!\Mux45~0_combout  & (\storeregister[21][18]~q )))) # (!temp_imemload_output_18 & (((\Mux45~0_combout ))))

	.dataa(\storeregister[21][18]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[29][18]~q ),
	.datad(\Mux45~0_combout ),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~1 .lut_mask = 16'hF388;
defparam \Mux45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N5
dffeas \storeregister[26][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][18] .is_wysiwyg = "true";
defparam \storeregister[26][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N4
cycloneive_lcell_comb \Mux45~3 (
// Equation(s):
// \Mux45~3_combout  = (\Mux45~2_combout  & (((\storeregister[30][18]~q )) # (!temp_imemload_output_19))) # (!\Mux45~2_combout  & (temp_imemload_output_19 & (\storeregister[26][18]~q )))

	.dataa(\Mux45~2_combout ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[26][18]~q ),
	.datad(\storeregister[30][18]~q ),
	.cin(gnd),
	.combout(\Mux45~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~3 .lut_mask = 16'hEA62;
defparam \Mux45~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N23
dffeas \storeregister[16][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][18] .is_wysiwyg = "true";
defparam \storeregister[16][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N22
cycloneive_lcell_comb \Mux45~4 (
// Equation(s):
// \Mux45~4_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[20][18]~q ))) # (!temp_imemload_output_18 & (\storeregister[16][18]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[16][18]~q ),
	.datad(\storeregister[20][18]~q ),
	.cin(gnd),
	.combout(\Mux45~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~4 .lut_mask = 16'hDC98;
defparam \Mux45~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N18
cycloneive_lcell_comb \Mux45~5 (
// Equation(s):
// \Mux45~5_combout  = (\Mux45~4_combout  & ((\storeregister[28][18]~q ) # ((!temp_imemload_output_19)))) # (!\Mux45~4_combout  & (((\storeregister[24][18]~q  & temp_imemload_output_19))))

	.dataa(\storeregister[28][18]~q ),
	.datab(\Mux45~4_combout ),
	.datac(\storeregister[24][18]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux45~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~5 .lut_mask = 16'hB8CC;
defparam \Mux45~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N26
cycloneive_lcell_comb \Mux45~6 (
// Equation(s):
// \Mux45~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\Mux45~3_combout )) # (!temp_imemload_output_17 & ((\Mux45~5_combout )))))

	.dataa(\Mux45~3_combout ),
	.datab(temp_imemload_output_16),
	.datac(\Mux45~5_combout ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux45~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~6 .lut_mask = 16'hEE30;
defparam \Mux45~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N12
cycloneive_lcell_comb \Mux45~12 (
// Equation(s):
// \Mux45~12_combout  = (temp_imemload_output_17 & ((\storeregister[10][18]~q ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((\storeregister[8][18]~q  & !temp_imemload_output_16))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[10][18]~q ),
	.datac(\storeregister[8][18]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux45~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~12 .lut_mask = 16'hAAD8;
defparam \Mux45~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N22
cycloneive_lcell_comb \Mux45~13 (
// Equation(s):
// \Mux45~13_combout  = (temp_imemload_output_16 & ((\Mux45~12_combout  & ((\storeregister[11][18]~q ))) # (!\Mux45~12_combout  & (\storeregister[9][18]~q )))) # (!temp_imemload_output_16 & (((\Mux45~12_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[9][18]~q ),
	.datac(\storeregister[11][18]~q ),
	.datad(\Mux45~12_combout ),
	.cin(gnd),
	.combout(\Mux45~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~13 .lut_mask = 16'hF588;
defparam \Mux45~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N0
cycloneive_lcell_comb \Mux45~15 (
// Equation(s):
// \Mux45~15_combout  = (\Mux45~14_combout ) # ((!temp_imemload_output_16 & (\storeregister[2][18]~q  & temp_imemload_output_17)))

	.dataa(\Mux45~14_combout ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[2][18]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux45~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~15 .lut_mask = 16'hBAAA;
defparam \Mux45~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N30
cycloneive_lcell_comb \Mux45~16 (
// Equation(s):
// \Mux45~16_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\Mux45~13_combout )) # (!temp_imemload_output_19 & ((\Mux45~15_combout )))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\Mux45~13_combout ),
	.datad(\Mux45~15_combout ),
	.cin(gnd),
	.combout(\Mux45~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~16 .lut_mask = 16'hD9C8;
defparam \Mux45~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N0
cycloneive_lcell_comb \Mux45~10 (
// Equation(s):
// \Mux45~10_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][18]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & ((\storeregister[4][18]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][18]~q ),
	.datad(\storeregister[4][18]~q ),
	.cin(gnd),
	.combout(\Mux45~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~10 .lut_mask = 16'hB9A8;
defparam \Mux45~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N10
cycloneive_lcell_comb \Mux45~11 (
// Equation(s):
// \Mux45~11_combout  = (\Mux45~10_combout  & (((\storeregister[7][18]~q )) # (!temp_imemload_output_17))) # (!\Mux45~10_combout  & (temp_imemload_output_17 & (\storeregister[6][18]~q )))

	.dataa(\Mux45~10_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[6][18]~q ),
	.datad(\storeregister[7][18]~q ),
	.cin(gnd),
	.combout(\Mux45~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~11 .lut_mask = 16'hEA62;
defparam \Mux45~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N10
cycloneive_lcell_comb \Mux45~17 (
// Equation(s):
// \Mux45~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][18]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][18]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[12][18]~q ),
	.datad(\storeregister[13][18]~q ),
	.cin(gnd),
	.combout(\Mux45~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~17 .lut_mask = 16'hDC98;
defparam \Mux45~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N16
cycloneive_lcell_comb \Mux45~18 (
// Equation(s):
// \Mux45~18_combout  = (\Mux45~17_combout  & ((\storeregister[15][18]~q ) # ((!temp_imemload_output_17)))) # (!\Mux45~17_combout  & (((\storeregister[14][18]~q  & temp_imemload_output_17))))

	.dataa(\storeregister[15][18]~q ),
	.datab(\storeregister[14][18]~q ),
	.datac(\Mux45~17_combout ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux45~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~18 .lut_mask = 16'hACF0;
defparam \Mux45~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N10
cycloneive_lcell_comb \Mux46~7 (
// Equation(s):
// \Mux46~7_combout  = (temp_imemload_output_18 & (((\storeregister[23][17]~q ) # (temp_imemload_output_19)))) # (!temp_imemload_output_18 & (\storeregister[19][17]~q  & ((!temp_imemload_output_19))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[19][17]~q ),
	.datac(\storeregister[23][17]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux46~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~7 .lut_mask = 16'hAAE4;
defparam \Mux46~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N12
cycloneive_lcell_comb \Mux46~8 (
// Equation(s):
// \Mux46~8_combout  = (\Mux46~7_combout  & (((\storeregister[31][17]~q ) # (!temp_imemload_output_19)))) # (!\Mux46~7_combout  & (\storeregister[27][17]~q  & ((temp_imemload_output_19))))

	.dataa(\storeregister[27][17]~q ),
	.datab(\Mux46~7_combout ),
	.datac(\storeregister[31][17]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux46~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~8 .lut_mask = 16'hE2CC;
defparam \Mux46~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N22
cycloneive_lcell_comb \Mux46~0 (
// Equation(s):
// \Mux46~0_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\storeregister[21][17]~q )) # (!temp_imemload_output_18 & ((\storeregister[17][17]~q )))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[21][17]~q ),
	.datad(\storeregister[17][17]~q ),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~0 .lut_mask = 16'hD9C8;
defparam \Mux46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N30
cycloneive_lcell_comb \Mux46~1 (
// Equation(s):
// \Mux46~1_combout  = (temp_imemload_output_19 & ((\Mux46~0_combout  & (\storeregister[29][17]~q )) # (!\Mux46~0_combout  & ((\storeregister[25][17]~q ))))) # (!temp_imemload_output_19 & (((\Mux46~0_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[29][17]~q ),
	.datac(\storeregister[25][17]~q ),
	.datad(\Mux46~0_combout ),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~1 .lut_mask = 16'hDDA0;
defparam \Mux46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N23
dffeas \storeregister[22][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][17] .is_wysiwyg = "true";
defparam \storeregister[22][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N18
cycloneive_lcell_comb \Mux46~3 (
// Equation(s):
// \Mux46~3_combout  = (\Mux46~2_combout  & (((\storeregister[30][17]~q ) # (!temp_imemload_output_18)))) # (!\Mux46~2_combout  & (\storeregister[22][17]~q  & ((temp_imemload_output_18))))

	.dataa(\Mux46~2_combout ),
	.datab(\storeregister[22][17]~q ),
	.datac(\storeregister[30][17]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux46~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~3 .lut_mask = 16'hE4AA;
defparam \Mux46~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N20
cycloneive_lcell_comb \storeregister[28][17]~feeder (
// Equation(s):
// \storeregister[28][17]~feeder_combout  = Mux14

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux14),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[28][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][17]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[28][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N21
dffeas \storeregister[28][17] (
	.clk(!CLK),
	.d(\storeregister[28][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][17] .is_wysiwyg = "true";
defparam \storeregister[28][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N8
cycloneive_lcell_comb \Mux46~4 (
// Equation(s):
// \Mux46~4_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[24][17]~q ))) # (!temp_imemload_output_19 & (\storeregister[16][17]~q ))))

	.dataa(\storeregister[16][17]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[24][17]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux46~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~4 .lut_mask = 16'hFC22;
defparam \Mux46~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N10
cycloneive_lcell_comb \Mux46~5 (
// Equation(s):
// \Mux46~5_combout  = (\Mux46~4_combout  & (((\storeregister[28][17]~q ) # (!temp_imemload_output_18)))) # (!\Mux46~4_combout  & (\storeregister[20][17]~q  & ((temp_imemload_output_18))))

	.dataa(\storeregister[20][17]~q ),
	.datab(\storeregister[28][17]~q ),
	.datac(\Mux46~4_combout ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux46~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~5 .lut_mask = 16'hCAF0;
defparam \Mux46~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N28
cycloneive_lcell_comb \Mux46~6 (
// Equation(s):
// \Mux46~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\Mux46~3_combout )) # (!temp_imemload_output_17 & ((\Mux46~5_combout )))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux46~3_combout ),
	.datac(temp_imemload_output_17),
	.datad(\Mux46~5_combout ),
	.cin(gnd),
	.combout(\Mux46~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~6 .lut_mask = 16'hE5E0;
defparam \Mux46~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N6
cycloneive_lcell_comb \Mux46~17 (
// Equation(s):
// \Mux46~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[13][17]~q )) # (!temp_imemload_output_16 & ((\storeregister[12][17]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[13][17]~q ),
	.datad(\storeregister[12][17]~q ),
	.cin(gnd),
	.combout(\Mux46~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~17 .lut_mask = 16'hD9C8;
defparam \Mux46~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N10
cycloneive_lcell_comb \Mux46~18 (
// Equation(s):
// \Mux46~18_combout  = (temp_imemload_output_17 & ((\Mux46~17_combout  & (\storeregister[15][17]~q )) # (!\Mux46~17_combout  & ((\storeregister[14][17]~q ))))) # (!temp_imemload_output_17 & (((\Mux46~17_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[15][17]~q ),
	.datac(\storeregister[14][17]~q ),
	.datad(\Mux46~17_combout ),
	.cin(gnd),
	.combout(\Mux46~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~18 .lut_mask = 16'hDDA0;
defparam \Mux46~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N30
cycloneive_lcell_comb \Mux46~14 (
// Equation(s):
// \Mux46~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][17]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][17]~q )))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[3][17]~q ),
	.datac(\storeregister[1][17]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux46~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~14 .lut_mask = 16'h88A0;
defparam \Mux46~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N16
cycloneive_lcell_comb \Mux46~15 (
// Equation(s):
// \Mux46~15_combout  = (\Mux46~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][17]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[2][17]~q ),
	.datac(\Mux46~14_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux46~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~15 .lut_mask = 16'hF0F8;
defparam \Mux46~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N6
cycloneive_lcell_comb \Mux46~12 (
// Equation(s):
// \Mux46~12_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][17]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & (\storeregister[4][17]~q )))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[4][17]~q ),
	.datad(\storeregister[5][17]~q ),
	.cin(gnd),
	.combout(\Mux46~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~12 .lut_mask = 16'hBA98;
defparam \Mux46~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N18
cycloneive_lcell_comb \Mux46~13 (
// Equation(s):
// \Mux46~13_combout  = (\Mux46~12_combout  & (((\storeregister[7][17]~q ) # (!temp_imemload_output_17)))) # (!\Mux46~12_combout  & (\storeregister[6][17]~q  & ((temp_imemload_output_17))))

	.dataa(\storeregister[6][17]~q ),
	.datab(\Mux46~12_combout ),
	.datac(\storeregister[7][17]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux46~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~13 .lut_mask = 16'hE2CC;
defparam \Mux46~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N12
cycloneive_lcell_comb \Mux46~16 (
// Equation(s):
// \Mux46~16_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19) # (\Mux46~13_combout )))) # (!temp_imemload_output_18 & (\Mux46~15_combout  & (!temp_imemload_output_19)))

	.dataa(\Mux46~15_combout ),
	.datab(temp_imemload_output_18),
	.datac(temp_imemload_output_19),
	.datad(\Mux46~13_combout ),
	.cin(gnd),
	.combout(\Mux46~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~16 .lut_mask = 16'hCEC2;
defparam \Mux46~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N28
cycloneive_lcell_comb \Mux46~10 (
// Equation(s):
// \Mux46~10_combout  = (temp_imemload_output_17 & (((\storeregister[10][17]~q ) # (temp_imemload_output_16)))) # (!temp_imemload_output_17 & (\storeregister[8][17]~q  & ((!temp_imemload_output_16))))

	.dataa(\storeregister[8][17]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[10][17]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux46~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~10 .lut_mask = 16'hCCE2;
defparam \Mux46~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N13
dffeas \storeregister[9][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][17] .is_wysiwyg = "true";
defparam \storeregister[9][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N12
cycloneive_lcell_comb \Mux46~11 (
// Equation(s):
// \Mux46~11_combout  = (temp_imemload_output_16 & ((\Mux46~10_combout  & ((\storeregister[11][17]~q ))) # (!\Mux46~10_combout  & (\storeregister[9][17]~q )))) # (!temp_imemload_output_16 & (\Mux46~10_combout ))

	.dataa(temp_imemload_output_16),
	.datab(\Mux46~10_combout ),
	.datac(\storeregister[9][17]~q ),
	.datad(\storeregister[11][17]~q ),
	.cin(gnd),
	.combout(\Mux46~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~11 .lut_mask = 16'hEC64;
defparam \Mux46~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N16
cycloneive_lcell_comb \Mux47~0 (
// Equation(s):
// \Mux47~0_combout  = (temp_imemload_output_19 & ((\storeregister[25][16]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\storeregister[17][16]~q  & !temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[25][16]~q ),
	.datac(\storeregister[17][16]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~0 .lut_mask = 16'hAAD8;
defparam \Mux47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N6
cycloneive_lcell_comb \Mux47~1 (
// Equation(s):
// \Mux47~1_combout  = (\Mux47~0_combout  & ((\storeregister[29][16]~q ) # ((!temp_imemload_output_18)))) # (!\Mux47~0_combout  & (((temp_imemload_output_18 & \storeregister[21][16]~q ))))

	.dataa(\Mux47~0_combout ),
	.datab(\storeregister[29][16]~q ),
	.datac(temp_imemload_output_18),
	.datad(\storeregister[21][16]~q ),
	.cin(gnd),
	.combout(\Mux47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~1 .lut_mask = 16'hDA8A;
defparam \Mux47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N31
dffeas \storeregister[19][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[19][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[19][16] .is_wysiwyg = "true";
defparam \storeregister[19][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N30
cycloneive_lcell_comb \Mux47~7 (
// Equation(s):
// \Mux47~7_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[27][16]~q ))) # (!temp_imemload_output_19 & (\storeregister[19][16]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[19][16]~q ),
	.datad(\storeregister[27][16]~q ),
	.cin(gnd),
	.combout(\Mux47~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~7 .lut_mask = 16'hDC98;
defparam \Mux47~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N18
cycloneive_lcell_comb \Mux47~8 (
// Equation(s):
// \Mux47~8_combout  = (temp_imemload_output_18 & ((\Mux47~7_combout  & ((\storeregister[31][16]~q ))) # (!\Mux47~7_combout  & (\storeregister[23][16]~q )))) # (!temp_imemload_output_18 & (((\Mux47~7_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[23][16]~q ),
	.datac(\storeregister[31][16]~q ),
	.datad(\Mux47~7_combout ),
	.cin(gnd),
	.combout(\Mux47~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~8 .lut_mask = 16'hF588;
defparam \Mux47~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N28
cycloneive_lcell_comb \storeregister[28][16]~feeder (
// Equation(s):
// \storeregister[28][16]~feeder_combout  = Mux15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux15),
	.cin(gnd),
	.combout(\storeregister[28][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][16]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[28][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N29
dffeas \storeregister[28][16] (
	.clk(!CLK),
	.d(\storeregister[28][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][16] .is_wysiwyg = "true";
defparam \storeregister[28][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N18
cycloneive_lcell_comb \Mux47~5 (
// Equation(s):
// \Mux47~5_combout  = (\Mux47~4_combout  & ((\storeregister[28][16]~q ) # ((!temp_imemload_output_19)))) # (!\Mux47~4_combout  & (((temp_imemload_output_19 & \storeregister[24][16]~q ))))

	.dataa(\Mux47~4_combout ),
	.datab(\storeregister[28][16]~q ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[24][16]~q ),
	.cin(gnd),
	.combout(\Mux47~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~5 .lut_mask = 16'hDA8A;
defparam \Mux47~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N24
cycloneive_lcell_comb \Mux47~2 (
// Equation(s):
// \Mux47~2_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\storeregister[22][16]~q )) # (!temp_imemload_output_18 & ((\storeregister[18][16]~q )))))

	.dataa(\storeregister[22][16]~q ),
	.datab(\storeregister[18][16]~q ),
	.datac(temp_imemload_output_19),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux47~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~2 .lut_mask = 16'hFA0C;
defparam \Mux47~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N12
cycloneive_lcell_comb \Mux47~3 (
// Equation(s):
// \Mux47~3_combout  = (temp_imemload_output_19 & ((\Mux47~2_combout  & ((\storeregister[30][16]~q ))) # (!\Mux47~2_combout  & (\storeregister[26][16]~q )))) # (!temp_imemload_output_19 & (((\Mux47~2_combout ))))

	.dataa(\storeregister[26][16]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[30][16]~q ),
	.datad(\Mux47~2_combout ),
	.cin(gnd),
	.combout(\Mux47~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~3 .lut_mask = 16'hF388;
defparam \Mux47~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N8
cycloneive_lcell_comb \Mux47~6 (
// Equation(s):
// \Mux47~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\Mux47~3_combout ))) # (!temp_imemload_output_17 & (\Mux47~5_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux47~5_combout ),
	.datac(temp_imemload_output_17),
	.datad(\Mux47~3_combout ),
	.cin(gnd),
	.combout(\Mux47~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~6 .lut_mask = 16'hF4A4;
defparam \Mux47~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N12
cycloneive_lcell_comb \Mux47~12 (
// Equation(s):
// \Mux47~12_combout  = (temp_imemload_output_17 & ((\storeregister[10][16]~q ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((!temp_imemload_output_16 & \storeregister[8][16]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[10][16]~q ),
	.datac(temp_imemload_output_16),
	.datad(\storeregister[8][16]~q ),
	.cin(gnd),
	.combout(\Mux47~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~12 .lut_mask = 16'hADA8;
defparam \Mux47~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N28
cycloneive_lcell_comb \Mux47~13 (
// Equation(s):
// \Mux47~13_combout  = (\Mux47~12_combout  & (((\storeregister[11][16]~q ) # (!temp_imemload_output_16)))) # (!\Mux47~12_combout  & (\storeregister[9][16]~q  & ((temp_imemload_output_16))))

	.dataa(\storeregister[9][16]~q ),
	.datab(\Mux47~12_combout ),
	.datac(\storeregister[11][16]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux47~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~13 .lut_mask = 16'hE2CC;
defparam \Mux47~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N0
cycloneive_lcell_comb \Mux47~14 (
// Equation(s):
// \Mux47~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][16]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][16]~q )))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[3][16]~q ),
	.datad(\storeregister[1][16]~q ),
	.cin(gnd),
	.combout(\Mux47~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~14 .lut_mask = 16'hA280;
defparam \Mux47~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N27
dffeas \storeregister[2][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][16] .is_wysiwyg = "true";
defparam \storeregister[2][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N26
cycloneive_lcell_comb \Mux47~15 (
// Equation(s):
// \Mux47~15_combout  = (\Mux47~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][16]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux47~14_combout ),
	.datac(\storeregister[2][16]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux47~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~15 .lut_mask = 16'hCCEC;
defparam \Mux47~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N28
cycloneive_lcell_comb \Mux47~16 (
// Equation(s):
// \Mux47~16_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\Mux47~13_combout )) # (!temp_imemload_output_19 & ((\Mux47~15_combout )))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\Mux47~13_combout ),
	.datad(\Mux47~15_combout ),
	.cin(gnd),
	.combout(\Mux47~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~16 .lut_mask = 16'hD9C8;
defparam \Mux47~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N24
cycloneive_lcell_comb \Mux47~10 (
// Equation(s):
// \Mux47~10_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[5][16]~q ))) # (!temp_imemload_output_16 & (\storeregister[4][16]~q ))))

	.dataa(\storeregister[4][16]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][16]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux47~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~10 .lut_mask = 16'hFC22;
defparam \Mux47~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N31
dffeas \storeregister[6][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][16] .is_wysiwyg = "true";
defparam \storeregister[6][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N30
cycloneive_lcell_comb \Mux47~11 (
// Equation(s):
// \Mux47~11_combout  = (\Mux47~10_combout  & (((\storeregister[7][16]~q )) # (!temp_imemload_output_17))) # (!\Mux47~10_combout  & (temp_imemload_output_17 & (\storeregister[6][16]~q )))

	.dataa(\Mux47~10_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[6][16]~q ),
	.datad(\storeregister[7][16]~q ),
	.cin(gnd),
	.combout(\Mux47~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~11 .lut_mask = 16'hEA62;
defparam \Mux47~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N18
cycloneive_lcell_comb \Mux47~17 (
// Equation(s):
// \Mux47~17_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[13][16]~q )) # (!temp_imemload_output_16 & ((\storeregister[12][16]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[13][16]~q ),
	.datac(\storeregister[12][16]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux47~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~17 .lut_mask = 16'hEE50;
defparam \Mux47~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N0
cycloneive_lcell_comb \Mux47~18 (
// Equation(s):
// \Mux47~18_combout  = (\Mux47~17_combout  & ((\storeregister[15][16]~q ) # ((!temp_imemload_output_17)))) # (!\Mux47~17_combout  & (((temp_imemload_output_17 & \storeregister[14][16]~q ))))

	.dataa(\storeregister[15][16]~q ),
	.datab(\Mux47~17_combout ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[14][16]~q ),
	.cin(gnd),
	.combout(\Mux47~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~18 .lut_mask = 16'hBC8C;
defparam \Mux47~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N31
dffeas \storeregister[17][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][31] .is_wysiwyg = "true";
defparam \storeregister[17][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N30
cycloneive_lcell_comb \Mux32~0 (
// Equation(s):
// \Mux32~0_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[21][31]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[17][31]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[17][31]~q ),
	.datad(\storeregister[21][31]~q ),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~0 .lut_mask = 16'hBA98;
defparam \Mux32~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N6
cycloneive_lcell_comb \Mux32~1 (
// Equation(s):
// \Mux32~1_combout  = (\Mux32~0_combout  & ((\storeregister[29][31]~q ) # ((!temp_imemload_output_19)))) # (!\Mux32~0_combout  & (((\storeregister[25][31]~q  & temp_imemload_output_19))))

	.dataa(\storeregister[29][31]~q ),
	.datab(\storeregister[25][31]~q ),
	.datac(\Mux32~0_combout ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~1 .lut_mask = 16'hACF0;
defparam \Mux32~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N6
cycloneive_lcell_comb \Mux32~7 (
// Equation(s):
// \Mux32~7_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[23][31]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[19][31]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[23][31]~q ),
	.datad(\storeregister[19][31]~q ),
	.cin(gnd),
	.combout(\Mux32~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~7 .lut_mask = 16'hB9A8;
defparam \Mux32~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N16
cycloneive_lcell_comb \Mux32~8 (
// Equation(s):
// \Mux32~8_combout  = (temp_imemload_output_19 & ((\Mux32~7_combout  & (\storeregister[31][31]~q )) # (!\Mux32~7_combout  & ((\storeregister[27][31]~q ))))) # (!temp_imemload_output_19 & (((\Mux32~7_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[31][31]~q ),
	.datac(\Mux32~7_combout ),
	.datad(\storeregister[27][31]~q ),
	.cin(gnd),
	.combout(\Mux32~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~8 .lut_mask = 16'hDAD0;
defparam \Mux32~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N30
cycloneive_lcell_comb \storeregister[16][31]~feeder (
// Equation(s):
// \storeregister[16][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux0),
	.cin(gnd),
	.combout(\storeregister[16][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[16][31]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[16][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N31
dffeas \storeregister[16][31] (
	.clk(!CLK),
	.d(\storeregister[16][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][31] .is_wysiwyg = "true";
defparam \storeregister[16][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N24
cycloneive_lcell_comb \Mux32~4 (
// Equation(s):
// \Mux32~4_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\storeregister[24][31]~q )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & (\storeregister[16][31]~q )))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[16][31]~q ),
	.datad(\storeregister[24][31]~q ),
	.cin(gnd),
	.combout(\Mux32~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~4 .lut_mask = 16'hBA98;
defparam \Mux32~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N26
cycloneive_lcell_comb \storeregister[28][31]~feeder (
// Equation(s):
// \storeregister[28][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux0),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[28][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][31]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[28][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N27
dffeas \storeregister[28][31] (
	.clk(!CLK),
	.d(\storeregister[28][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][31] .is_wysiwyg = "true";
defparam \storeregister[28][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N12
cycloneive_lcell_comb \Mux32~5 (
// Equation(s):
// \Mux32~5_combout  = (temp_imemload_output_18 & ((\Mux32~4_combout  & (\storeregister[28][31]~q )) # (!\Mux32~4_combout  & ((\storeregister[20][31]~q ))))) # (!temp_imemload_output_18 & (\Mux32~4_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux32~4_combout ),
	.datac(\storeregister[28][31]~q ),
	.datad(\storeregister[20][31]~q ),
	.cin(gnd),
	.combout(\Mux32~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~5 .lut_mask = 16'hE6C4;
defparam \Mux32~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N14
cycloneive_lcell_comb \storeregister[22][31]~feeder (
// Equation(s):
// \storeregister[22][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux0),
	.cin(gnd),
	.combout(\storeregister[22][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[22][31]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[22][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N15
dffeas \storeregister[22][31] (
	.clk(!CLK),
	.d(\storeregister[22][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][31] .is_wysiwyg = "true";
defparam \storeregister[22][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N14
cycloneive_lcell_comb \Mux32~3 (
// Equation(s):
// \Mux32~3_combout  = (\Mux32~2_combout  & (((\storeregister[30][31]~q )) # (!temp_imemload_output_18))) # (!\Mux32~2_combout  & (temp_imemload_output_18 & (\storeregister[22][31]~q )))

	.dataa(\Mux32~2_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[22][31]~q ),
	.datad(\storeregister[30][31]~q ),
	.cin(gnd),
	.combout(\Mux32~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~3 .lut_mask = 16'hEA62;
defparam \Mux32~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N26
cycloneive_lcell_comb \Mux32~6 (
// Equation(s):
// \Mux32~6_combout  = (temp_imemload_output_17 & (((\Mux32~3_combout ) # (temp_imemload_output_16)))) # (!temp_imemload_output_17 & (\Mux32~5_combout  & ((!temp_imemload_output_16))))

	.dataa(\Mux32~5_combout ),
	.datab(\Mux32~3_combout ),
	.datac(temp_imemload_output_17),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux32~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~6 .lut_mask = 16'hF0CA;
defparam \Mux32~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N17
dffeas \storeregister[10][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][31] .is_wysiwyg = "true";
defparam \storeregister[10][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N16
cycloneive_lcell_comb \Mux32~10 (
// Equation(s):
// \Mux32~10_combout  = (temp_imemload_output_17 & (((\storeregister[10][31]~q ) # (temp_imemload_output_16)))) # (!temp_imemload_output_17 & (\storeregister[8][31]~q  & ((!temp_imemload_output_16))))

	.dataa(\storeregister[8][31]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[10][31]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux32~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~10 .lut_mask = 16'hCCE2;
defparam \Mux32~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N16
cycloneive_lcell_comb \Mux32~11 (
// Equation(s):
// \Mux32~11_combout  = (temp_imemload_output_16 & ((\Mux32~10_combout  & (\storeregister[11][31]~q )) # (!\Mux32~10_combout  & ((\storeregister[9][31]~q ))))) # (!temp_imemload_output_16 & (((\Mux32~10_combout ))))

	.dataa(\storeregister[11][31]~q ),
	.datab(temp_imemload_output_16),
	.datac(\Mux32~10_combout ),
	.datad(\storeregister[9][31]~q ),
	.cin(gnd),
	.combout(\Mux32~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~11 .lut_mask = 16'hBCB0;
defparam \Mux32~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N14
cycloneive_lcell_comb \storeregister[13][31]~feeder (
// Equation(s):
// \storeregister[13][31]~feeder_combout  = Mux0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux0),
	.cin(gnd),
	.combout(\storeregister[13][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[13][31]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[13][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N15
dffeas \storeregister[13][31] (
	.clk(!CLK),
	.d(\storeregister[13][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[13][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[13][31] .is_wysiwyg = "true";
defparam \storeregister[13][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N24
cycloneive_lcell_comb \Mux32~17 (
// Equation(s):
// \Mux32~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][31]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][31]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[12][31]~q ),
	.datad(\storeregister[13][31]~q ),
	.cin(gnd),
	.combout(\Mux32~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~17 .lut_mask = 16'hDC98;
defparam \Mux32~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N4
cycloneive_lcell_comb \Mux32~18 (
// Equation(s):
// \Mux32~18_combout  = (temp_imemload_output_17 & ((\Mux32~17_combout  & ((\storeregister[15][31]~q ))) # (!\Mux32~17_combout  & (\storeregister[14][31]~q )))) # (!temp_imemload_output_17 & (((\Mux32~17_combout ))))

	.dataa(\storeregister[14][31]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[15][31]~q ),
	.datad(\Mux32~17_combout ),
	.cin(gnd),
	.combout(\Mux32~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~18 .lut_mask = 16'hF388;
defparam \Mux32~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N18
cycloneive_lcell_comb \Mux32~12 (
// Equation(s):
// \Mux32~12_combout  = (temp_imemload_output_16 & ((\storeregister[5][31]~q ) # ((temp_imemload_output_17)))) # (!temp_imemload_output_16 & (((\storeregister[4][31]~q  & !temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[5][31]~q ),
	.datac(\storeregister[4][31]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux32~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~12 .lut_mask = 16'hAAD8;
defparam \Mux32~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N16
cycloneive_lcell_comb \Mux32~13 (
// Equation(s):
// \Mux32~13_combout  = (temp_imemload_output_17 & ((\Mux32~12_combout  & (\storeregister[7][31]~q )) # (!\Mux32~12_combout  & ((\storeregister[6][31]~q ))))) # (!temp_imemload_output_17 & (\Mux32~12_combout ))

	.dataa(temp_imemload_output_17),
	.datab(\Mux32~12_combout ),
	.datac(\storeregister[7][31]~q ),
	.datad(\storeregister[6][31]~q ),
	.cin(gnd),
	.combout(\Mux32~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~13 .lut_mask = 16'hE6C4;
defparam \Mux32~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N20
cycloneive_lcell_comb \Mux32~15 (
// Equation(s):
// \Mux32~15_combout  = (\Mux32~14_combout ) # ((\storeregister[2][31]~q  & (temp_imemload_output_17 & !temp_imemload_output_16)))

	.dataa(\Mux32~14_combout ),
	.datab(\storeregister[2][31]~q ),
	.datac(temp_imemload_output_17),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux32~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~15 .lut_mask = 16'hAAEA;
defparam \Mux32~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N14
cycloneive_lcell_comb \Mux32~16 (
// Equation(s):
// \Mux32~16_combout  = (temp_imemload_output_18 & ((\Mux32~13_combout ) # ((temp_imemload_output_19)))) # (!temp_imemload_output_18 & (((\Mux32~15_combout  & !temp_imemload_output_19))))

	.dataa(\Mux32~13_combout ),
	.datab(\Mux32~15_combout ),
	.datac(temp_imemload_output_18),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux32~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~16 .lut_mask = 16'hF0AC;
defparam \Mux32~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N12
cycloneive_lcell_comb \Mux33~0 (
// Equation(s):
// \Mux33~0_combout  = (temp_imemload_output_19 & (((\storeregister[25][30]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[17][30]~q  & ((!temp_imemload_output_18))))

	.dataa(\storeregister[17][30]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[25][30]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~0 .lut_mask = 16'hCCE2;
defparam \Mux33~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N2
cycloneive_lcell_comb \Mux33~1 (
// Equation(s):
// \Mux33~1_combout  = (\Mux33~0_combout  & (((\storeregister[29][30]~q ) # (!temp_imemload_output_18)))) # (!\Mux33~0_combout  & (\storeregister[21][30]~q  & ((temp_imemload_output_18))))

	.dataa(\Mux33~0_combout ),
	.datab(\storeregister[21][30]~q ),
	.datac(\storeregister[29][30]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~1 .lut_mask = 16'hE4AA;
defparam \Mux33~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N2
cycloneive_lcell_comb \Mux33~4 (
// Equation(s):
// \Mux33~4_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[20][30]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[16][30]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[20][30]~q ),
	.datad(\storeregister[16][30]~q ),
	.cin(gnd),
	.combout(\Mux33~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~4 .lut_mask = 16'hB9A8;
defparam \Mux33~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N10
cycloneive_lcell_comb \Mux33~5 (
// Equation(s):
// \Mux33~5_combout  = (temp_imemload_output_19 & ((\Mux33~4_combout  & (\storeregister[28][30]~q )) # (!\Mux33~4_combout  & ((\storeregister[24][30]~q ))))) # (!temp_imemload_output_19 & (((\Mux33~4_combout ))))

	.dataa(\storeregister[28][30]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[24][30]~q ),
	.datad(\Mux33~4_combout ),
	.cin(gnd),
	.combout(\Mux33~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~5 .lut_mask = 16'hBBC0;
defparam \Mux33~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N31
dffeas \storeregister[18][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][30] .is_wysiwyg = "true";
defparam \storeregister[18][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N12
cycloneive_lcell_comb \storeregister[22][30]~feeder (
// Equation(s):
// \storeregister[22][30]~feeder_combout  = Mux1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux1),
	.cin(gnd),
	.combout(\storeregister[22][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[22][30]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[22][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N13
dffeas \storeregister[22][30] (
	.clk(!CLK),
	.d(\storeregister[22][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][30] .is_wysiwyg = "true";
defparam \storeregister[22][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N30
cycloneive_lcell_comb \Mux33~2 (
// Equation(s):
// \Mux33~2_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[22][30]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[18][30]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[18][30]~q ),
	.datad(\storeregister[22][30]~q ),
	.cin(gnd),
	.combout(\Mux33~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~2 .lut_mask = 16'hBA98;
defparam \Mux33~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N18
cycloneive_lcell_comb \Mux33~3 (
// Equation(s):
// \Mux33~3_combout  = (temp_imemload_output_19 & ((\Mux33~2_combout  & ((\storeregister[30][30]~q ))) # (!\Mux33~2_combout  & (\storeregister[26][30]~q )))) # (!temp_imemload_output_19 & (((\Mux33~2_combout ))))

	.dataa(\storeregister[26][30]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[30][30]~q ),
	.datad(\Mux33~2_combout ),
	.cin(gnd),
	.combout(\Mux33~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~3 .lut_mask = 16'hF388;
defparam \Mux33~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N28
cycloneive_lcell_comb \Mux33~6 (
// Equation(s):
// \Mux33~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\Mux33~3_combout ))) # (!temp_imemload_output_17 & (\Mux33~5_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux33~5_combout ),
	.datac(\Mux33~3_combout ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux33~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~6 .lut_mask = 16'hFA44;
defparam \Mux33~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N26
cycloneive_lcell_comb \Mux33~7 (
// Equation(s):
// \Mux33~7_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\storeregister[27][30]~q )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & ((\storeregister[19][30]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[27][30]~q ),
	.datad(\storeregister[19][30]~q ),
	.cin(gnd),
	.combout(\Mux33~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~7 .lut_mask = 16'hB9A8;
defparam \Mux33~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N24
cycloneive_lcell_comb \Mux33~8 (
// Equation(s):
// \Mux33~8_combout  = (\Mux33~7_combout  & (((\storeregister[31][30]~q )) # (!temp_imemload_output_18))) # (!\Mux33~7_combout  & (temp_imemload_output_18 & (\storeregister[23][30]~q )))

	.dataa(\Mux33~7_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[23][30]~q ),
	.datad(\storeregister[31][30]~q ),
	.cin(gnd),
	.combout(\Mux33~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~8 .lut_mask = 16'hEA62;
defparam \Mux33~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y40_N17
dffeas \storeregister[5][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][30] .is_wysiwyg = "true";
defparam \storeregister[5][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N16
cycloneive_lcell_comb \Mux33~10 (
// Equation(s):
// \Mux33~10_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[5][30]~q ))) # (!temp_imemload_output_16 & (\storeregister[4][30]~q ))))

	.dataa(\storeregister[4][30]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][30]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux33~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~10 .lut_mask = 16'hFC22;
defparam \Mux33~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N2
cycloneive_lcell_comb \Mux33~11 (
// Equation(s):
// \Mux33~11_combout  = (temp_imemload_output_17 & ((\Mux33~10_combout  & (\storeregister[7][30]~q )) # (!\Mux33~10_combout  & ((\storeregister[6][30]~q ))))) # (!temp_imemload_output_17 & (((\Mux33~10_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[7][30]~q ),
	.datac(\storeregister[6][30]~q ),
	.datad(\Mux33~10_combout ),
	.cin(gnd),
	.combout(\Mux33~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~11 .lut_mask = 16'hDDA0;
defparam \Mux33~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N10
cycloneive_lcell_comb \Mux33~17 (
// Equation(s):
// \Mux33~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[13][30]~q )) # (!temp_imemload_output_16 & ((\storeregister[12][30]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[13][30]~q ),
	.datad(\storeregister[12][30]~q ),
	.cin(gnd),
	.combout(\Mux33~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~17 .lut_mask = 16'hD9C8;
defparam \Mux33~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N8
cycloneive_lcell_comb \Mux33~18 (
// Equation(s):
// \Mux33~18_combout  = (\Mux33~17_combout  & (((\storeregister[15][30]~q ) # (!temp_imemload_output_17)))) # (!\Mux33~17_combout  & (\storeregister[14][30]~q  & ((temp_imemload_output_17))))

	.dataa(\Mux33~17_combout ),
	.datab(\storeregister[14][30]~q ),
	.datac(\storeregister[15][30]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux33~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~18 .lut_mask = 16'hE4AA;
defparam \Mux33~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y40_N5
dffeas \storeregister[8][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][30] .is_wysiwyg = "true";
defparam \storeregister[8][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N4
cycloneive_lcell_comb \Mux33~12 (
// Equation(s):
// \Mux33~12_combout  = (temp_imemload_output_17 & ((temp_imemload_output_16) # ((\storeregister[10][30]~q )))) # (!temp_imemload_output_17 & (!temp_imemload_output_16 & (\storeregister[8][30]~q )))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[8][30]~q ),
	.datad(\storeregister[10][30]~q ),
	.cin(gnd),
	.combout(\Mux33~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~12 .lut_mask = 16'hBA98;
defparam \Mux33~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N28
cycloneive_lcell_comb \Mux33~13 (
// Equation(s):
// \Mux33~13_combout  = (\Mux33~12_combout  & (((\storeregister[11][30]~q ) # (!temp_imemload_output_16)))) # (!\Mux33~12_combout  & (\storeregister[9][30]~q  & ((temp_imemload_output_16))))

	.dataa(\storeregister[9][30]~q ),
	.datab(\Mux33~12_combout ),
	.datac(\storeregister[11][30]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux33~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~13 .lut_mask = 16'hE2CC;
defparam \Mux33~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N14
cycloneive_lcell_comb \Mux33~14 (
// Equation(s):
// \Mux33~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][30]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][30]~q )))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[3][30]~q ),
	.datac(\storeregister[1][30]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux33~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~14 .lut_mask = 16'h88A0;
defparam \Mux33~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N10
cycloneive_lcell_comb \Mux33~15 (
// Equation(s):
// \Mux33~15_combout  = (\Mux33~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][30]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[2][30]~q ),
	.datac(\Mux33~14_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux33~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~15 .lut_mask = 16'hF0F8;
defparam \Mux33~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N12
cycloneive_lcell_comb \Mux33~16 (
// Equation(s):
// \Mux33~16_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\Mux33~13_combout )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & ((\Mux33~15_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\Mux33~13_combout ),
	.datad(\Mux33~15_combout ),
	.cin(gnd),
	.combout(\Mux33~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~16 .lut_mask = 16'hB9A8;
defparam \Mux33~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N26
cycloneive_lcell_comb \Mux34~7 (
// Equation(s):
// \Mux34~7_combout  = (temp_imemload_output_18 & (((\storeregister[23][29]~q ) # (temp_imemload_output_19)))) # (!temp_imemload_output_18 & (\storeregister[19][29]~q  & ((!temp_imemload_output_19))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[19][29]~q ),
	.datac(\storeregister[23][29]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux34~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~7 .lut_mask = 16'hAAE4;
defparam \Mux34~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N14
cycloneive_lcell_comb \Mux34~8 (
// Equation(s):
// \Mux34~8_combout  = (temp_imemload_output_19 & ((\Mux34~7_combout  & (\storeregister[31][29]~q )) # (!\Mux34~7_combout  & ((\storeregister[27][29]~q ))))) # (!temp_imemload_output_19 & (((\Mux34~7_combout ))))

	.dataa(\storeregister[31][29]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[27][29]~q ),
	.datad(\Mux34~7_combout ),
	.cin(gnd),
	.combout(\Mux34~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~8 .lut_mask = 16'hBBC0;
defparam \Mux34~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N18
cycloneive_lcell_comb \Mux34~3 (
// Equation(s):
// \Mux34~3_combout  = (\Mux34~2_combout  & (((\storeregister[30][29]~q )) # (!temp_imemload_output_18))) # (!\Mux34~2_combout  & (temp_imemload_output_18 & ((\storeregister[22][29]~q ))))

	.dataa(\Mux34~2_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[30][29]~q ),
	.datad(\storeregister[22][29]~q ),
	.cin(gnd),
	.combout(\Mux34~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~3 .lut_mask = 16'hE6A2;
defparam \Mux34~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N26
cycloneive_lcell_comb \storeregister[28][29]~feeder (
// Equation(s):
// \storeregister[28][29]~feeder_combout  = Mux2

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux2),
	.cin(gnd),
	.combout(\storeregister[28][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[28][29]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[28][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N27
dffeas \storeregister[28][29] (
	.clk(!CLK),
	.d(\storeregister[28][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[28][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[28][29] .is_wysiwyg = "true";
defparam \storeregister[28][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N0
cycloneive_lcell_comb \storeregister[20][29]~feeder (
// Equation(s):
// \storeregister[20][29]~feeder_combout  = Mux2

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux2),
	.cin(gnd),
	.combout(\storeregister[20][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][29]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[20][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N1
dffeas \storeregister[20][29] (
	.clk(!CLK),
	.d(\storeregister[20][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][29] .is_wysiwyg = "true";
defparam \storeregister[20][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N6
cycloneive_lcell_comb \Mux34~5 (
// Equation(s):
// \Mux34~5_combout  = (\Mux34~4_combout  & (((\storeregister[28][29]~q )) # (!temp_imemload_output_18))) # (!\Mux34~4_combout  & (temp_imemload_output_18 & ((\storeregister[20][29]~q ))))

	.dataa(\Mux34~4_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[28][29]~q ),
	.datad(\storeregister[20][29]~q ),
	.cin(gnd),
	.combout(\Mux34~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~5 .lut_mask = 16'hE6A2;
defparam \Mux34~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N18
cycloneive_lcell_comb \Mux34~6 (
// Equation(s):
// \Mux34~6_combout  = (temp_imemload_output_17 & ((\Mux34~3_combout ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((!temp_imemload_output_16 & \Mux34~5_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\Mux34~3_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux34~5_combout ),
	.cin(gnd),
	.combout(\Mux34~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~6 .lut_mask = 16'hADA8;
defparam \Mux34~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N10
cycloneive_lcell_comb \Mux34~0 (
// Equation(s):
// \Mux34~0_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[21][29]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[17][29]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[17][29]~q ),
	.datad(\storeregister[21][29]~q ),
	.cin(gnd),
	.combout(\Mux34~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~0 .lut_mask = 16'hBA98;
defparam \Mux34~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N28
cycloneive_lcell_comb \Mux34~1 (
// Equation(s):
// \Mux34~1_combout  = (temp_imemload_output_19 & ((\Mux34~0_combout  & ((\storeregister[29][29]~q ))) # (!\Mux34~0_combout  & (\storeregister[25][29]~q )))) # (!temp_imemload_output_19 & (((\Mux34~0_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[25][29]~q ),
	.datac(\Mux34~0_combout ),
	.datad(\storeregister[29][29]~q ),
	.cin(gnd),
	.combout(\Mux34~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~1 .lut_mask = 16'hF858;
defparam \Mux34~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N8
cycloneive_lcell_comb \Mux34~10 (
// Equation(s):
// \Mux34~10_combout  = (temp_imemload_output_17 & (((\storeregister[10][29]~q ) # (temp_imemload_output_16)))) # (!temp_imemload_output_17 & (\storeregister[8][29]~q  & ((!temp_imemload_output_16))))

	.dataa(\storeregister[8][29]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[10][29]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux34~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~10 .lut_mask = 16'hCCE2;
defparam \Mux34~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N20
cycloneive_lcell_comb \Mux34~11 (
// Equation(s):
// \Mux34~11_combout  = (temp_imemload_output_16 & ((\Mux34~10_combout  & ((\storeregister[11][29]~q ))) # (!\Mux34~10_combout  & (\storeregister[9][29]~q )))) # (!temp_imemload_output_16 & (((\Mux34~10_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[9][29]~q ),
	.datac(\storeregister[11][29]~q ),
	.datad(\Mux34~10_combout ),
	.cin(gnd),
	.combout(\Mux34~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~11 .lut_mask = 16'hF588;
defparam \Mux34~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N22
cycloneive_lcell_comb \Mux34~13 (
// Equation(s):
// \Mux34~13_combout  = (\Mux34~12_combout  & (((\storeregister[7][29]~q )) # (!temp_imemload_output_17))) # (!\Mux34~12_combout  & (temp_imemload_output_17 & ((\storeregister[6][29]~q ))))

	.dataa(\Mux34~12_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[7][29]~q ),
	.datad(\storeregister[6][29]~q ),
	.cin(gnd),
	.combout(\Mux34~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~13 .lut_mask = 16'hE6A2;
defparam \Mux34~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N21
dffeas \storeregister[3][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][29] .is_wysiwyg = "true";
defparam \storeregister[3][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N23
dffeas \storeregister[1][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][29] .is_wysiwyg = "true";
defparam \storeregister[1][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N22
cycloneive_lcell_comb \Mux34~14 (
// Equation(s):
// \Mux34~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][29]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][29]~q )))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[3][29]~q ),
	.datac(\storeregister[1][29]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux34~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~14 .lut_mask = 16'h88A0;
defparam \Mux34~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N10
cycloneive_lcell_comb \Mux34~15 (
// Equation(s):
// \Mux34~15_combout  = (\Mux34~14_combout ) # ((temp_imemload_output_17 & (!temp_imemload_output_16 & \storeregister[2][29]~q )))

	.dataa(temp_imemload_output_17),
	.datab(\Mux34~14_combout ),
	.datac(temp_imemload_output_16),
	.datad(\storeregister[2][29]~q ),
	.cin(gnd),
	.combout(\Mux34~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~15 .lut_mask = 16'hCECC;
defparam \Mux34~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N8
cycloneive_lcell_comb \Mux34~16 (
// Equation(s):
// \Mux34~16_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\Mux34~13_combout )) # (!temp_imemload_output_18 & ((\Mux34~15_combout )))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\Mux34~13_combout ),
	.datad(\Mux34~15_combout ),
	.cin(gnd),
	.combout(\Mux34~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~16 .lut_mask = 16'hD9C8;
defparam \Mux34~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N28
cycloneive_lcell_comb \Mux34~17 (
// Equation(s):
// \Mux34~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[13][29]~q )) # (!temp_imemload_output_16 & ((\storeregister[12][29]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[13][29]~q ),
	.datad(\storeregister[12][29]~q ),
	.cin(gnd),
	.combout(\Mux34~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~17 .lut_mask = 16'hD9C8;
defparam \Mux34~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N30
cycloneive_lcell_comb \Mux34~18 (
// Equation(s):
// \Mux34~18_combout  = (\Mux34~17_combout  & (((\storeregister[15][29]~q )) # (!temp_imemload_output_17))) # (!\Mux34~17_combout  & (temp_imemload_output_17 & (\storeregister[14][29]~q )))

	.dataa(\Mux34~17_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[14][29]~q ),
	.datad(\storeregister[15][29]~q ),
	.cin(gnd),
	.combout(\Mux34~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~18 .lut_mask = 16'hEA62;
defparam \Mux34~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N2
cycloneive_lcell_comb \Mux35~7 (
// Equation(s):
// \Mux35~7_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[27][28]~q ))) # (!temp_imemload_output_19 & (\storeregister[19][28]~q ))))

	.dataa(\storeregister[19][28]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[27][28]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux35~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~7 .lut_mask = 16'hFC22;
defparam \Mux35~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N8
cycloneive_lcell_comb \Mux35~8 (
// Equation(s):
// \Mux35~8_combout  = (temp_imemload_output_18 & ((\Mux35~7_combout  & ((\storeregister[31][28]~q ))) # (!\Mux35~7_combout  & (\storeregister[23][28]~q )))) # (!temp_imemload_output_18 & (((\Mux35~7_combout ))))

	.dataa(\storeregister[23][28]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[31][28]~q ),
	.datad(\Mux35~7_combout ),
	.cin(gnd),
	.combout(\Mux35~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~8 .lut_mask = 16'hF388;
defparam \Mux35~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N11
dffeas \storeregister[18][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][28] .is_wysiwyg = "true";
defparam \storeregister[18][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N4
cycloneive_lcell_comb \storeregister[22][28]~feeder (
// Equation(s):
// \storeregister[22][28]~feeder_combout  = Mux3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux3),
	.cin(gnd),
	.combout(\storeregister[22][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[22][28]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[22][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N5
dffeas \storeregister[22][28] (
	.clk(!CLK),
	.d(\storeregister[22][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][28] .is_wysiwyg = "true";
defparam \storeregister[22][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N10
cycloneive_lcell_comb \Mux35~2 (
// Equation(s):
// \Mux35~2_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[22][28]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[18][28]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[18][28]~q ),
	.datad(\storeregister[22][28]~q ),
	.cin(gnd),
	.combout(\Mux35~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~2 .lut_mask = 16'hBA98;
defparam \Mux35~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N16
cycloneive_lcell_comb \Mux35~3 (
// Equation(s):
// \Mux35~3_combout  = (temp_imemload_output_19 & ((\Mux35~2_combout  & (\storeregister[30][28]~q )) # (!\Mux35~2_combout  & ((\storeregister[26][28]~q ))))) # (!temp_imemload_output_19 & (((\Mux35~2_combout ))))

	.dataa(\storeregister[30][28]~q ),
	.datab(\storeregister[26][28]~q ),
	.datac(temp_imemload_output_19),
	.datad(\Mux35~2_combout ),
	.cin(gnd),
	.combout(\Mux35~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~3 .lut_mask = 16'hAFC0;
defparam \Mux35~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N10
cycloneive_lcell_comb \Mux35~4 (
// Equation(s):
// \Mux35~4_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[20][28]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[16][28]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[20][28]~q ),
	.datad(\storeregister[16][28]~q ),
	.cin(gnd),
	.combout(\Mux35~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~4 .lut_mask = 16'hB9A8;
defparam \Mux35~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N16
cycloneive_lcell_comb \Mux35~5 (
// Equation(s):
// \Mux35~5_combout  = (\Mux35~4_combout  & ((\storeregister[28][28]~q ) # ((!temp_imemload_output_19)))) # (!\Mux35~4_combout  & (((temp_imemload_output_19 & \storeregister[24][28]~q ))))

	.dataa(\storeregister[28][28]~q ),
	.datab(\Mux35~4_combout ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[24][28]~q ),
	.cin(gnd),
	.combout(\Mux35~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~5 .lut_mask = 16'hBC8C;
defparam \Mux35~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N30
cycloneive_lcell_comb \Mux35~6 (
// Equation(s):
// \Mux35~6_combout  = (temp_imemload_output_16 & (temp_imemload_output_17)) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\Mux35~3_combout )) # (!temp_imemload_output_17 & ((\Mux35~5_combout )))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\Mux35~3_combout ),
	.datad(\Mux35~5_combout ),
	.cin(gnd),
	.combout(\Mux35~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~6 .lut_mask = 16'hD9C8;
defparam \Mux35~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N8
cycloneive_lcell_comb \Mux35~0 (
// Equation(s):
// \Mux35~0_combout  = (temp_imemload_output_19 & (((\storeregister[25][28]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[17][28]~q  & ((!temp_imemload_output_18))))

	.dataa(\storeregister[17][28]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[25][28]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux35~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~0 .lut_mask = 16'hCCE2;
defparam \Mux35~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N4
cycloneive_lcell_comb \Mux35~1 (
// Equation(s):
// \Mux35~1_combout  = (\Mux35~0_combout  & (((\storeregister[29][28]~q ) # (!temp_imemload_output_18)))) # (!\Mux35~0_combout  & (\storeregister[21][28]~q  & (temp_imemload_output_18)))

	.dataa(\Mux35~0_combout ),
	.datab(\storeregister[21][28]~q ),
	.datac(temp_imemload_output_18),
	.datad(\storeregister[29][28]~q ),
	.cin(gnd),
	.combout(\Mux35~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~1 .lut_mask = 16'hEA4A;
defparam \Mux35~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y41_N21
dffeas \storeregister[5][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][28] .is_wysiwyg = "true";
defparam \storeregister[5][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N20
cycloneive_lcell_comb \Mux35~10 (
// Equation(s):
// \Mux35~10_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[5][28]~q ))) # (!temp_imemload_output_16 & (\storeregister[4][28]~q ))))

	.dataa(\storeregister[4][28]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][28]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux35~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~10 .lut_mask = 16'hFC22;
defparam \Mux35~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N24
cycloneive_lcell_comb \Mux35~11 (
// Equation(s):
// \Mux35~11_combout  = (temp_imemload_output_17 & ((\Mux35~10_combout  & (\storeregister[7][28]~q )) # (!\Mux35~10_combout  & ((\storeregister[6][28]~q ))))) # (!temp_imemload_output_17 & (((\Mux35~10_combout ))))

	.dataa(\storeregister[7][28]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[6][28]~q ),
	.datad(\Mux35~10_combout ),
	.cin(gnd),
	.combout(\Mux35~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~11 .lut_mask = 16'hBBC0;
defparam \Mux35~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N7
dffeas \storeregister[1][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][28] .is_wysiwyg = "true";
defparam \storeregister[1][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N6
cycloneive_lcell_comb \Mux35~14 (
// Equation(s):
// \Mux35~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[3][28]~q ))) # (!temp_imemload_output_17 & (\storeregister[1][28]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[1][28]~q ),
	.datad(\storeregister[3][28]~q ),
	.cin(gnd),
	.combout(\Mux35~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~14 .lut_mask = 16'hC840;
defparam \Mux35~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N6
cycloneive_lcell_comb \Mux35~15 (
// Equation(s):
// \Mux35~15_combout  = (\Mux35~14_combout ) # ((!temp_imemload_output_16 & (temp_imemload_output_17 & \storeregister[2][28]~q )))

	.dataa(temp_imemload_output_16),
	.datab(\Mux35~14_combout ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[2][28]~q ),
	.cin(gnd),
	.combout(\Mux35~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~15 .lut_mask = 16'hDCCC;
defparam \Mux35~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N10
cycloneive_lcell_comb \Mux35~13 (
// Equation(s):
// \Mux35~13_combout  = (\Mux35~12_combout  & (((\storeregister[11][28]~q ) # (!temp_imemload_output_16)))) # (!\Mux35~12_combout  & (\storeregister[9][28]~q  & ((temp_imemload_output_16))))

	.dataa(\Mux35~12_combout ),
	.datab(\storeregister[9][28]~q ),
	.datac(\storeregister[11][28]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux35~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~13 .lut_mask = 16'hE4AA;
defparam \Mux35~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N22
cycloneive_lcell_comb \Mux35~16 (
// Equation(s):
// \Mux35~16_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\Mux35~13_combout ))) # (!temp_imemload_output_19 & (\Mux35~15_combout ))))

	.dataa(\Mux35~15_combout ),
	.datab(temp_imemload_output_18),
	.datac(temp_imemload_output_19),
	.datad(\Mux35~13_combout ),
	.cin(gnd),
	.combout(\Mux35~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~16 .lut_mask = 16'hF2C2;
defparam \Mux35~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y40_N28
cycloneive_lcell_comb \Mux35~17 (
// Equation(s):
// \Mux35~17_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][28]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][28]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[12][28]~q ),
	.datac(temp_imemload_output_16),
	.datad(\storeregister[13][28]~q ),
	.cin(gnd),
	.combout(\Mux35~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~17 .lut_mask = 16'hF4A4;
defparam \Mux35~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y40_N14
cycloneive_lcell_comb \Mux35~18 (
// Equation(s):
// \Mux35~18_combout  = (\Mux35~17_combout  & ((\storeregister[15][28]~q ) # ((!temp_imemload_output_17)))) # (!\Mux35~17_combout  & (((temp_imemload_output_17 & \storeregister[14][28]~q ))))

	.dataa(\storeregister[15][28]~q ),
	.datab(\Mux35~17_combout ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[14][28]~q ),
	.cin(gnd),
	.combout(\Mux35~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~18 .lut_mask = 16'hBC8C;
defparam \Mux35~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N21
dffeas \storeregister[17][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][26] .is_wysiwyg = "true";
defparam \storeregister[17][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N20
cycloneive_lcell_comb \Mux37~0 (
// Equation(s):
// \Mux37~0_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[25][26]~q ))) # (!temp_imemload_output_19 & (\storeregister[17][26]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[17][26]~q ),
	.datad(\storeregister[25][26]~q ),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~0 .lut_mask = 16'hDC98;
defparam \Mux37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N26
cycloneive_lcell_comb \Mux37~1 (
// Equation(s):
// \Mux37~1_combout  = (temp_imemload_output_18 & ((\Mux37~0_combout  & ((\storeregister[29][26]~q ))) # (!\Mux37~0_combout  & (\storeregister[21][26]~q )))) # (!temp_imemload_output_18 & (((\Mux37~0_combout ))))

	.dataa(\storeregister[21][26]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[29][26]~q ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\Mux37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~1 .lut_mask = 16'hF388;
defparam \Mux37~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N27
dffeas \storeregister[18][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][26] .is_wysiwyg = "true";
defparam \storeregister[18][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N26
cycloneive_lcell_comb \Mux37~2 (
// Equation(s):
// \Mux37~2_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[22][26]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[18][26]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[18][26]~q ),
	.datad(\storeregister[22][26]~q ),
	.cin(gnd),
	.combout(\Mux37~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~2 .lut_mask = 16'hBA98;
defparam \Mux37~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N22
cycloneive_lcell_comb \Mux37~3 (
// Equation(s):
// \Mux37~3_combout  = (temp_imemload_output_19 & ((\Mux37~2_combout  & ((\storeregister[30][26]~q ))) # (!\Mux37~2_combout  & (\storeregister[26][26]~q )))) # (!temp_imemload_output_19 & (((\Mux37~2_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[26][26]~q ),
	.datac(\Mux37~2_combout ),
	.datad(\storeregister[30][26]~q ),
	.cin(gnd),
	.combout(\Mux37~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~3 .lut_mask = 16'hF858;
defparam \Mux37~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N19
dffeas \storeregister[20][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][26] .is_wysiwyg = "true";
defparam \storeregister[20][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N18
cycloneive_lcell_comb \Mux37~4 (
// Equation(s):
// \Mux37~4_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[20][26]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[16][26]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[20][26]~q ),
	.datad(\storeregister[16][26]~q ),
	.cin(gnd),
	.combout(\Mux37~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~4 .lut_mask = 16'hB9A8;
defparam \Mux37~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N18
cycloneive_lcell_comb \Mux37~5 (
// Equation(s):
// \Mux37~5_combout  = (temp_imemload_output_19 & ((\Mux37~4_combout  & ((\storeregister[28][26]~q ))) # (!\Mux37~4_combout  & (\storeregister[24][26]~q )))) # (!temp_imemload_output_19 & (\Mux37~4_combout ))

	.dataa(temp_imemload_output_19),
	.datab(\Mux37~4_combout ),
	.datac(\storeregister[24][26]~q ),
	.datad(\storeregister[28][26]~q ),
	.cin(gnd),
	.combout(\Mux37~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~5 .lut_mask = 16'hEC64;
defparam \Mux37~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N14
cycloneive_lcell_comb \Mux37~6 (
// Equation(s):
// \Mux37~6_combout  = (temp_imemload_output_17 & ((\Mux37~3_combout ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((!temp_imemload_output_16 & \Mux37~5_combout ))))

	.dataa(\Mux37~3_combout ),
	.datab(temp_imemload_output_17),
	.datac(temp_imemload_output_16),
	.datad(\Mux37~5_combout ),
	.cin(gnd),
	.combout(\Mux37~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~6 .lut_mask = 16'hCBC8;
defparam \Mux37~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N24
cycloneive_lcell_comb \Mux37~7 (
// Equation(s):
// \Mux37~7_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[27][26]~q ))) # (!temp_imemload_output_19 & (\storeregister[19][26]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[19][26]~q ),
	.datac(\storeregister[27][26]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux37~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~7 .lut_mask = 16'hFA44;
defparam \Mux37~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N2
cycloneive_lcell_comb \Mux37~8 (
// Equation(s):
// \Mux37~8_combout  = (temp_imemload_output_18 & ((\Mux37~7_combout  & (\storeregister[31][26]~q )) # (!\Mux37~7_combout  & ((\storeregister[23][26]~q ))))) # (!temp_imemload_output_18 & (((\Mux37~7_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[31][26]~q ),
	.datac(\Mux37~7_combout ),
	.datad(\storeregister[23][26]~q ),
	.cin(gnd),
	.combout(\Mux37~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~8 .lut_mask = 16'hDAD0;
defparam \Mux37~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N15
dffeas \storeregister[1][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][26] .is_wysiwyg = "true";
defparam \storeregister[1][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N14
cycloneive_lcell_comb \Mux37~14 (
// Equation(s):
// \Mux37~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][26]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][26]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[3][26]~q ),
	.datac(\storeregister[1][26]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux37~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~14 .lut_mask = 16'hD800;
defparam \Mux37~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N12
cycloneive_lcell_comb \Mux37~15 (
// Equation(s):
// \Mux37~15_combout  = (\Mux37~14_combout ) # ((temp_imemload_output_17 & (!temp_imemload_output_16 & \storeregister[2][26]~q )))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[2][26]~q ),
	.datad(\Mux37~14_combout ),
	.cin(gnd),
	.combout(\Mux37~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~15 .lut_mask = 16'hFF20;
defparam \Mux37~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N5
dffeas \storeregister[8][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][26] .is_wysiwyg = "true";
defparam \storeregister[8][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N4
cycloneive_lcell_comb \Mux37~12 (
// Equation(s):
// \Mux37~12_combout  = (temp_imemload_output_17 & ((\storeregister[10][26]~q ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((\storeregister[8][26]~q  & !temp_imemload_output_16))))

	.dataa(\storeregister[10][26]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[8][26]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux37~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~12 .lut_mask = 16'hCCB8;
defparam \Mux37~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N22
cycloneive_lcell_comb \Mux37~13 (
// Equation(s):
// \Mux37~13_combout  = (temp_imemload_output_16 & ((\Mux37~12_combout  & ((\storeregister[11][26]~q ))) # (!\Mux37~12_combout  & (\storeregister[9][26]~q )))) # (!temp_imemload_output_16 & (((\Mux37~12_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[9][26]~q ),
	.datac(\storeregister[11][26]~q ),
	.datad(\Mux37~12_combout ),
	.cin(gnd),
	.combout(\Mux37~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~13 .lut_mask = 16'hF588;
defparam \Mux37~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N6
cycloneive_lcell_comb \Mux37~16 (
// Equation(s):
// \Mux37~16_combout  = (temp_imemload_output_19 & (((\Mux37~13_combout ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\Mux37~15_combout  & ((!temp_imemload_output_18))))

	.dataa(\Mux37~15_combout ),
	.datab(temp_imemload_output_19),
	.datac(\Mux37~13_combout ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux37~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~16 .lut_mask = 16'hCCE2;
defparam \Mux37~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y41_N29
dffeas \storeregister[5][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][26] .is_wysiwyg = "true";
defparam \storeregister[5][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y41_N3
dffeas \storeregister[4][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][26] .is_wysiwyg = "true";
defparam \storeregister[4][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N28
cycloneive_lcell_comb \Mux37~10 (
// Equation(s):
// \Mux37~10_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][26]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & ((\storeregister[4][26]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][26]~q ),
	.datad(\storeregister[4][26]~q ),
	.cin(gnd),
	.combout(\Mux37~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~10 .lut_mask = 16'hB9A8;
defparam \Mux37~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N0
cycloneive_lcell_comb \Mux37~11 (
// Equation(s):
// \Mux37~11_combout  = (\Mux37~10_combout  & ((\storeregister[7][26]~q ) # ((!temp_imemload_output_17)))) # (!\Mux37~10_combout  & (((\storeregister[6][26]~q  & temp_imemload_output_17))))

	.dataa(\storeregister[7][26]~q ),
	.datab(\Mux37~10_combout ),
	.datac(\storeregister[6][26]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux37~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~11 .lut_mask = 16'hB8CC;
defparam \Mux37~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N0
cycloneive_lcell_comb \Mux37~17 (
// Equation(s):
// \Mux37~17_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][26]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][26]~q ))))

	.dataa(\storeregister[12][26]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[13][26]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux37~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~17 .lut_mask = 16'hFC22;
defparam \Mux37~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N10
cycloneive_lcell_comb \Mux37~18 (
// Equation(s):
// \Mux37~18_combout  = (\Mux37~17_combout  & (((\storeregister[15][26]~q )) # (!temp_imemload_output_17))) # (!\Mux37~17_combout  & (temp_imemload_output_17 & (\storeregister[14][26]~q )))

	.dataa(\Mux37~17_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[14][26]~q ),
	.datad(\storeregister[15][26]~q ),
	.cin(gnd),
	.combout(\Mux37~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~18 .lut_mask = 16'hEA62;
defparam \Mux37~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N10
cycloneive_lcell_comb \Mux38~7 (
// Equation(s):
// \Mux38~7_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\storeregister[23][25]~q )) # (!temp_imemload_output_18 & ((\storeregister[19][25]~q )))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[23][25]~q ),
	.datad(\storeregister[19][25]~q ),
	.cin(gnd),
	.combout(\Mux38~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~7 .lut_mask = 16'hD9C8;
defparam \Mux38~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N8
cycloneive_lcell_comb \Mux38~8 (
// Equation(s):
// \Mux38~8_combout  = (\Mux38~7_combout  & (((\storeregister[31][25]~q ) # (!temp_imemload_output_19)))) # (!\Mux38~7_combout  & (\storeregister[27][25]~q  & ((temp_imemload_output_19))))

	.dataa(\Mux38~7_combout ),
	.datab(\storeregister[27][25]~q ),
	.datac(\storeregister[31][25]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux38~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~8 .lut_mask = 16'hE4AA;
defparam \Mux38~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N10
cycloneive_lcell_comb \Mux38~0 (
// Equation(s):
// \Mux38~0_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[21][25]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[17][25]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[17][25]~q ),
	.datad(\storeregister[21][25]~q ),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~0 .lut_mask = 16'hBA98;
defparam \Mux38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N0
cycloneive_lcell_comb \Mux38~1 (
// Equation(s):
// \Mux38~1_combout  = (\Mux38~0_combout  & (((\storeregister[29][25]~q )) # (!temp_imemload_output_19))) # (!\Mux38~0_combout  & (temp_imemload_output_19 & ((\storeregister[25][25]~q ))))

	.dataa(\Mux38~0_combout ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[29][25]~q ),
	.datad(\storeregister[25][25]~q ),
	.cin(gnd),
	.combout(\Mux38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~1 .lut_mask = 16'hE6A2;
defparam \Mux38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N4
cycloneive_lcell_comb \Mux38~3 (
// Equation(s):
// \Mux38~3_combout  = (\Mux38~2_combout  & (((\storeregister[30][25]~q )) # (!temp_imemload_output_18))) # (!\Mux38~2_combout  & (temp_imemload_output_18 & (\storeregister[22][25]~q )))

	.dataa(\Mux38~2_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[22][25]~q ),
	.datad(\storeregister[30][25]~q ),
	.cin(gnd),
	.combout(\Mux38~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~3 .lut_mask = 16'hEA62;
defparam \Mux38~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N17
dffeas \storeregister[24][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][25] .is_wysiwyg = "true";
defparam \storeregister[24][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N16
cycloneive_lcell_comb \Mux38~4 (
// Equation(s):
// \Mux38~4_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[24][25]~q ))) # (!temp_imemload_output_19 & (\storeregister[16][25]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[16][25]~q ),
	.datac(\storeregister[24][25]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux38~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~4 .lut_mask = 16'hFA44;
defparam \Mux38~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N30
cycloneive_lcell_comb \Mux38~5 (
// Equation(s):
// \Mux38~5_combout  = (temp_imemload_output_18 & ((\Mux38~4_combout  & (\storeregister[28][25]~q )) # (!\Mux38~4_combout  & ((\storeregister[20][25]~q ))))) # (!temp_imemload_output_18 & (((\Mux38~4_combout ))))

	.dataa(\storeregister[28][25]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[20][25]~q ),
	.datad(\Mux38~4_combout ),
	.cin(gnd),
	.combout(\Mux38~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~5 .lut_mask = 16'hBBC0;
defparam \Mux38~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N16
cycloneive_lcell_comb \Mux38~6 (
// Equation(s):
// \Mux38~6_combout  = (temp_imemload_output_17 & ((temp_imemload_output_16) # ((\Mux38~3_combout )))) # (!temp_imemload_output_17 & (!temp_imemload_output_16 & ((\Mux38~5_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\Mux38~3_combout ),
	.datad(\Mux38~5_combout ),
	.cin(gnd),
	.combout(\Mux38~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~6 .lut_mask = 16'hB9A8;
defparam \Mux38~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N6
cycloneive_lcell_comb \Mux38~13 (
// Equation(s):
// \Mux38~13_combout  = (\Mux38~12_combout  & (((\storeregister[7][25]~q )) # (!temp_imemload_output_17))) # (!\Mux38~12_combout  & (temp_imemload_output_17 & ((\storeregister[6][25]~q ))))

	.dataa(\Mux38~12_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[7][25]~q ),
	.datad(\storeregister[6][25]~q ),
	.cin(gnd),
	.combout(\Mux38~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~13 .lut_mask = 16'hE6A2;
defparam \Mux38~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N23
dffeas \storeregister[1][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][25] .is_wysiwyg = "true";
defparam \storeregister[1][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N22
cycloneive_lcell_comb \Mux38~14 (
// Equation(s):
// \Mux38~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][25]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][25]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[3][25]~q ),
	.datac(\storeregister[1][25]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux38~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~14 .lut_mask = 16'hD800;
defparam \Mux38~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N20
cycloneive_lcell_comb \Mux38~15 (
// Equation(s):
// \Mux38~15_combout  = (\Mux38~14_combout ) # ((!temp_imemload_output_16 & (temp_imemload_output_17 & \storeregister[2][25]~q )))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\Mux38~14_combout ),
	.datad(\storeregister[2][25]~q ),
	.cin(gnd),
	.combout(\Mux38~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~15 .lut_mask = 16'hF4F0;
defparam \Mux38~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N26
cycloneive_lcell_comb \Mux38~16 (
// Equation(s):
// \Mux38~16_combout  = (temp_imemload_output_18 & ((\Mux38~13_combout ) # ((temp_imemload_output_19)))) # (!temp_imemload_output_18 & (((!temp_imemload_output_19 & \Mux38~15_combout ))))

	.dataa(\Mux38~13_combout ),
	.datab(temp_imemload_output_18),
	.datac(temp_imemload_output_19),
	.datad(\Mux38~15_combout ),
	.cin(gnd),
	.combout(\Mux38~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~16 .lut_mask = 16'hCBC8;
defparam \Mux38~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N24
cycloneive_lcell_comb \Mux38~17 (
// Equation(s):
// \Mux38~17_combout  = (temp_imemload_output_16 & (((\storeregister[13][25]~q ) # (temp_imemload_output_17)))) # (!temp_imemload_output_16 & (\storeregister[12][25]~q  & ((!temp_imemload_output_17))))

	.dataa(\storeregister[12][25]~q ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[13][25]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux38~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~17 .lut_mask = 16'hCCE2;
defparam \Mux38~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N0
cycloneive_lcell_comb \Mux38~18 (
// Equation(s):
// \Mux38~18_combout  = (\Mux38~17_combout  & ((\storeregister[15][25]~q ) # ((!temp_imemload_output_17)))) # (!\Mux38~17_combout  & (((\storeregister[14][25]~q  & temp_imemload_output_17))))

	.dataa(\storeregister[15][25]~q ),
	.datab(\Mux38~17_combout ),
	.datac(\storeregister[14][25]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux38~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~18 .lut_mask = 16'hB8CC;
defparam \Mux38~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N15
dffeas \storeregister[10][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][25] .is_wysiwyg = "true";
defparam \storeregister[10][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N14
cycloneive_lcell_comb \Mux38~10 (
// Equation(s):
// \Mux38~10_combout  = (temp_imemload_output_17 & (((\storeregister[10][25]~q ) # (temp_imemload_output_16)))) # (!temp_imemload_output_17 & (\storeregister[8][25]~q  & ((!temp_imemload_output_16))))

	.dataa(\storeregister[8][25]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[10][25]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux38~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~10 .lut_mask = 16'hCCE2;
defparam \Mux38~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N28
cycloneive_lcell_comb \Mux38~11 (
// Equation(s):
// \Mux38~11_combout  = (\Mux38~10_combout  & (((\storeregister[11][25]~q )) # (!temp_imemload_output_16))) # (!\Mux38~10_combout  & (temp_imemload_output_16 & (\storeregister[9][25]~q )))

	.dataa(\Mux38~10_combout ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[9][25]~q ),
	.datad(\storeregister[11][25]~q ),
	.cin(gnd),
	.combout(\Mux38~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~11 .lut_mask = 16'hEA62;
defparam \Mux38~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N0
cycloneive_lcell_comb \storeregister[20][24]~feeder (
// Equation(s):
// \storeregister[20][24]~feeder_combout  = Mux7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux7),
	.cin(gnd),
	.combout(\storeregister[20][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][24]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[20][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N1
dffeas \storeregister[20][24] (
	.clk(!CLK),
	.d(\storeregister[20][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][24] .is_wysiwyg = "true";
defparam \storeregister[20][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N14
cycloneive_lcell_comb \Mux39~4 (
// Equation(s):
// \Mux39~4_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[20][24]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[16][24]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[16][24]~q ),
	.datad(\storeregister[20][24]~q ),
	.cin(gnd),
	.combout(\Mux39~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~4 .lut_mask = 16'hBA98;
defparam \Mux39~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N2
cycloneive_lcell_comb \Mux39~5 (
// Equation(s):
// \Mux39~5_combout  = (temp_imemload_output_19 & ((\Mux39~4_combout  & (\storeregister[28][24]~q )) # (!\Mux39~4_combout  & ((\storeregister[24][24]~q ))))) # (!temp_imemload_output_19 & (((\Mux39~4_combout ))))

	.dataa(\storeregister[28][24]~q ),
	.datab(\storeregister[24][24]~q ),
	.datac(temp_imemload_output_19),
	.datad(\Mux39~4_combout ),
	.cin(gnd),
	.combout(\Mux39~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~5 .lut_mask = 16'hAFC0;
defparam \Mux39~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N8
cycloneive_lcell_comb \Mux39~3 (
// Equation(s):
// \Mux39~3_combout  = (\Mux39~2_combout  & (((\storeregister[30][24]~q )) # (!temp_imemload_output_19))) # (!\Mux39~2_combout  & (temp_imemload_output_19 & (\storeregister[26][24]~q )))

	.dataa(\Mux39~2_combout ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[26][24]~q ),
	.datad(\storeregister[30][24]~q ),
	.cin(gnd),
	.combout(\Mux39~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~3 .lut_mask = 16'hEA62;
defparam \Mux39~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N12
cycloneive_lcell_comb \Mux39~6 (
// Equation(s):
// \Mux39~6_combout  = (temp_imemload_output_17 & (((\Mux39~3_combout ) # (temp_imemload_output_16)))) # (!temp_imemload_output_17 & (\Mux39~5_combout  & ((!temp_imemload_output_16))))

	.dataa(temp_imemload_output_17),
	.datab(\Mux39~5_combout ),
	.datac(\Mux39~3_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux39~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~6 .lut_mask = 16'hAAE4;
defparam \Mux39~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N29
dffeas \storeregister[17][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][24] .is_wysiwyg = "true";
defparam \storeregister[17][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N28
cycloneive_lcell_comb \Mux39~0 (
// Equation(s):
// \Mux39~0_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[25][24]~q ))) # (!temp_imemload_output_19 & (\storeregister[17][24]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[17][24]~q ),
	.datad(\storeregister[25][24]~q ),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~0 .lut_mask = 16'hDC98;
defparam \Mux39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N0
cycloneive_lcell_comb \Mux39~1 (
// Equation(s):
// \Mux39~1_combout  = (\Mux39~0_combout  & (((\storeregister[29][24]~q ) # (!temp_imemload_output_18)))) # (!\Mux39~0_combout  & (\storeregister[21][24]~q  & ((temp_imemload_output_18))))

	.dataa(\storeregister[21][24]~q ),
	.datab(\Mux39~0_combout ),
	.datac(\storeregister[29][24]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~1 .lut_mask = 16'hE2CC;
defparam \Mux39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N6
cycloneive_lcell_comb \storeregister[23][24]~feeder (
// Equation(s):
// \storeregister[23][24]~feeder_combout  = Mux7

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux7),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[23][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][24]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[23][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N7
dffeas \storeregister[23][24] (
	.clk(!CLK),
	.d(\storeregister[23][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][24] .is_wysiwyg = "true";
defparam \storeregister[23][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N24
cycloneive_lcell_comb \Mux39~7 (
// Equation(s):
// \Mux39~7_combout  = (temp_imemload_output_19 & (((\storeregister[27][24]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[19][24]~q  & ((!temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[19][24]~q ),
	.datac(\storeregister[27][24]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux39~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~7 .lut_mask = 16'hAAE4;
defparam \Mux39~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N16
cycloneive_lcell_comb \Mux39~8 (
// Equation(s):
// \Mux39~8_combout  = (temp_imemload_output_18 & ((\Mux39~7_combout  & (\storeregister[31][24]~q )) # (!\Mux39~7_combout  & ((\storeregister[23][24]~q ))))) # (!temp_imemload_output_18 & (((\Mux39~7_combout ))))

	.dataa(\storeregister[31][24]~q ),
	.datab(\storeregister[23][24]~q ),
	.datac(temp_imemload_output_18),
	.datad(\Mux39~7_combout ),
	.cin(gnd),
	.combout(\Mux39~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~8 .lut_mask = 16'hAFC0;
defparam \Mux39~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y41_N13
dffeas \storeregister[5][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][24] .is_wysiwyg = "true";
defparam \storeregister[5][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N12
cycloneive_lcell_comb \Mux39~10 (
// Equation(s):
// \Mux39~10_combout  = (temp_imemload_output_16 & (((\storeregister[5][24]~q ) # (temp_imemload_output_17)))) # (!temp_imemload_output_16 & (\storeregister[4][24]~q  & ((!temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[4][24]~q ),
	.datac(\storeregister[5][24]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux39~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~10 .lut_mask = 16'hAAE4;
defparam \Mux39~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y41_N27
dffeas \storeregister[6][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][24] .is_wysiwyg = "true";
defparam \storeregister[6][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N26
cycloneive_lcell_comb \Mux39~11 (
// Equation(s):
// \Mux39~11_combout  = (\Mux39~10_combout  & ((\storeregister[7][24]~q ) # ((!temp_imemload_output_17)))) # (!\Mux39~10_combout  & (((\storeregister[6][24]~q  & temp_imemload_output_17))))

	.dataa(\Mux39~10_combout ),
	.datab(\storeregister[7][24]~q ),
	.datac(\storeregister[6][24]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux39~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~11 .lut_mask = 16'hD8AA;
defparam \Mux39~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N15
dffeas \storeregister[12][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[12][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[12][24] .is_wysiwyg = "true";
defparam \storeregister[12][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N14
cycloneive_lcell_comb \Mux39~17 (
// Equation(s):
// \Mux39~17_combout  = (temp_imemload_output_16 & ((\storeregister[13][24]~q ) # ((temp_imemload_output_17)))) # (!temp_imemload_output_16 & (((\storeregister[12][24]~q  & !temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[13][24]~q ),
	.datac(\storeregister[12][24]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux39~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~17 .lut_mask = 16'hAAD8;
defparam \Mux39~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N30
cycloneive_lcell_comb \Mux39~18 (
// Equation(s):
// \Mux39~18_combout  = (\Mux39~17_combout  & (((\storeregister[15][24]~q ) # (!temp_imemload_output_17)))) # (!\Mux39~17_combout  & (\storeregister[14][24]~q  & (temp_imemload_output_17)))

	.dataa(\Mux39~17_combout ),
	.datab(\storeregister[14][24]~q ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[15][24]~q ),
	.cin(gnd),
	.combout(\Mux39~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~18 .lut_mask = 16'hEA4A;
defparam \Mux39~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N20
cycloneive_lcell_comb \Mux39~12 (
// Equation(s):
// \Mux39~12_combout  = (temp_imemload_output_16 & (temp_imemload_output_17)) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[10][24]~q ))) # (!temp_imemload_output_17 & (\storeregister[8][24]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[8][24]~q ),
	.datad(\storeregister[10][24]~q ),
	.cin(gnd),
	.combout(\Mux39~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~12 .lut_mask = 16'hDC98;
defparam \Mux39~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N30
cycloneive_lcell_comb \Mux39~13 (
// Equation(s):
// \Mux39~13_combout  = (temp_imemload_output_16 & ((\Mux39~12_combout  & ((\storeregister[11][24]~q ))) # (!\Mux39~12_combout  & (\storeregister[9][24]~q )))) # (!temp_imemload_output_16 & (((\Mux39~12_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[9][24]~q ),
	.datac(\storeregister[11][24]~q ),
	.datad(\Mux39~12_combout ),
	.cin(gnd),
	.combout(\Mux39~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~13 .lut_mask = 16'hF588;
defparam \Mux39~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N11
dffeas \storeregister[1][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][24] .is_wysiwyg = "true";
defparam \storeregister[1][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N10
cycloneive_lcell_comb \Mux39~14 (
// Equation(s):
// \Mux39~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][24]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][24]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[3][24]~q ),
	.datac(\storeregister[1][24]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux39~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~14 .lut_mask = 16'hD800;
defparam \Mux39~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N10
cycloneive_lcell_comb \Mux39~15 (
// Equation(s):
// \Mux39~15_combout  = (\Mux39~14_combout ) # ((!temp_imemload_output_16 & (temp_imemload_output_17 & \storeregister[2][24]~q )))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\Mux39~14_combout ),
	.datad(\storeregister[2][24]~q ),
	.cin(gnd),
	.combout(\Mux39~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~15 .lut_mask = 16'hF4F0;
defparam \Mux39~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N12
cycloneive_lcell_comb \Mux39~16 (
// Equation(s):
// \Mux39~16_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\Mux39~13_combout )) # (!temp_imemload_output_19 & ((\Mux39~15_combout )))))

	.dataa(\Mux39~13_combout ),
	.datab(temp_imemload_output_18),
	.datac(temp_imemload_output_19),
	.datad(\Mux39~15_combout ),
	.cin(gnd),
	.combout(\Mux39~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~16 .lut_mask = 16'hE3E0;
defparam \Mux39~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N8
cycloneive_lcell_comb \Mux40~4 (
// Equation(s):
// \Mux40~4_combout  = (temp_imemload_output_19 & (((\storeregister[24][23]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[16][23]~q  & ((!temp_imemload_output_18))))

	.dataa(\storeregister[16][23]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[24][23]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux40~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~4 .lut_mask = 16'hCCE2;
defparam \Mux40~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N20
cycloneive_lcell_comb \Mux40~5 (
// Equation(s):
// \Mux40~5_combout  = (temp_imemload_output_18 & ((\Mux40~4_combout  & (\storeregister[28][23]~q )) # (!\Mux40~4_combout  & ((\storeregister[20][23]~q ))))) # (!temp_imemload_output_18 & (((\Mux40~4_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[28][23]~q ),
	.datac(\storeregister[20][23]~q ),
	.datad(\Mux40~4_combout ),
	.cin(gnd),
	.combout(\Mux40~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~5 .lut_mask = 16'hDDA0;
defparam \Mux40~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N23
dffeas \storeregister[22][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][23] .is_wysiwyg = "true";
defparam \storeregister[22][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N3
dffeas \storeregister[18][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][23] .is_wysiwyg = "true";
defparam \storeregister[18][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N28
cycloneive_lcell_comb \Mux40~2 (
// Equation(s):
// \Mux40~2_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[26][23]~q ))) # (!temp_imemload_output_19 & (\storeregister[18][23]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[18][23]~q ),
	.datac(\storeregister[26][23]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux40~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~2 .lut_mask = 16'hFA44;
defparam \Mux40~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N22
cycloneive_lcell_comb \Mux40~3 (
// Equation(s):
// \Mux40~3_combout  = (temp_imemload_output_18 & ((\Mux40~2_combout  & (\storeregister[30][23]~q )) # (!\Mux40~2_combout  & ((\storeregister[22][23]~q ))))) # (!temp_imemload_output_18 & (((\Mux40~2_combout ))))

	.dataa(\storeregister[30][23]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[22][23]~q ),
	.datad(\Mux40~2_combout ),
	.cin(gnd),
	.combout(\Mux40~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~3 .lut_mask = 16'hBBC0;
defparam \Mux40~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N18
cycloneive_lcell_comb \Mux40~6 (
// Equation(s):
// \Mux40~6_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16) # (\Mux40~3_combout )))) # (!temp_imemload_output_17 & (\Mux40~5_combout  & (!temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux40~5_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux40~3_combout ),
	.cin(gnd),
	.combout(\Mux40~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~6 .lut_mask = 16'hAEA4;
defparam \Mux40~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N28
cycloneive_lcell_comb \Mux40~7 (
// Equation(s):
// \Mux40~7_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[23][23]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[19][23]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[23][23]~q ),
	.datad(\storeregister[19][23]~q ),
	.cin(gnd),
	.combout(\Mux40~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~7 .lut_mask = 16'hB9A8;
defparam \Mux40~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N16
cycloneive_lcell_comb \Mux40~8 (
// Equation(s):
// \Mux40~8_combout  = (temp_imemload_output_19 & ((\Mux40~7_combout  & (\storeregister[31][23]~q )) # (!\Mux40~7_combout  & ((\storeregister[27][23]~q ))))) # (!temp_imemload_output_19 & (\Mux40~7_combout ))

	.dataa(temp_imemload_output_19),
	.datab(\Mux40~7_combout ),
	.datac(\storeregister[31][23]~q ),
	.datad(\storeregister[27][23]~q ),
	.cin(gnd),
	.combout(\Mux40~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~8 .lut_mask = 16'hE6C4;
defparam \Mux40~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N6
cycloneive_lcell_comb \Mux40~0 (
// Equation(s):
// \Mux40~0_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[21][23]~q ))) # (!temp_imemload_output_18 & (\storeregister[17][23]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[17][23]~q ),
	.datad(\storeregister[21][23]~q ),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~0 .lut_mask = 16'hDC98;
defparam \Mux40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N4
cycloneive_lcell_comb \Mux40~1 (
// Equation(s):
// \Mux40~1_combout  = (temp_imemload_output_19 & ((\Mux40~0_combout  & (\storeregister[29][23]~q )) # (!\Mux40~0_combout  & ((\storeregister[25][23]~q ))))) # (!temp_imemload_output_19 & (((\Mux40~0_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[29][23]~q ),
	.datac(\storeregister[25][23]~q ),
	.datad(\Mux40~0_combout ),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~1 .lut_mask = 16'hDDA0;
defparam \Mux40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N6
cycloneive_lcell_comb \Mux40~17 (
// Equation(s):
// \Mux40~17_combout  = (temp_imemload_output_16 & ((\storeregister[13][23]~q ) # ((temp_imemload_output_17)))) # (!temp_imemload_output_16 & (((\storeregister[12][23]~q  & !temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[13][23]~q ),
	.datac(\storeregister[12][23]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux40~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~17 .lut_mask = 16'hAAD8;
defparam \Mux40~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N18
cycloneive_lcell_comb \Mux40~18 (
// Equation(s):
// \Mux40~18_combout  = (temp_imemload_output_17 & ((\Mux40~17_combout  & ((\storeregister[15][23]~q ))) # (!\Mux40~17_combout  & (\storeregister[14][23]~q )))) # (!temp_imemload_output_17 & (\Mux40~17_combout ))

	.dataa(temp_imemload_output_17),
	.datab(\Mux40~17_combout ),
	.datac(\storeregister[14][23]~q ),
	.datad(\storeregister[15][23]~q ),
	.cin(gnd),
	.combout(\Mux40~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~18 .lut_mask = 16'hEC64;
defparam \Mux40~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N14
cycloneive_lcell_comb \Mux40~13 (
// Equation(s):
// \Mux40~13_combout  = (\Mux40~12_combout  & (((\storeregister[7][23]~q ) # (!temp_imemload_output_17)))) # (!\Mux40~12_combout  & (\storeregister[6][23]~q  & ((temp_imemload_output_17))))

	.dataa(\Mux40~12_combout ),
	.datab(\storeregister[6][23]~q ),
	.datac(\storeregister[7][23]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux40~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~13 .lut_mask = 16'hE4AA;
defparam \Mux40~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N18
cycloneive_lcell_comb \Mux40~14 (
// Equation(s):
// \Mux40~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][23]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][23]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[3][23]~q ),
	.datac(\storeregister[1][23]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux40~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~14 .lut_mask = 16'hD800;
defparam \Mux40~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N10
cycloneive_lcell_comb \Mux40~15 (
// Equation(s):
// \Mux40~15_combout  = (\Mux40~14_combout ) # ((!temp_imemload_output_16 & (\storeregister[2][23]~q  & temp_imemload_output_17)))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[2][23]~q ),
	.datac(temp_imemload_output_17),
	.datad(\Mux40~14_combout ),
	.cin(gnd),
	.combout(\Mux40~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~15 .lut_mask = 16'hFF40;
defparam \Mux40~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N4
cycloneive_lcell_comb \Mux40~16 (
// Equation(s):
// \Mux40~16_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\Mux40~13_combout )) # (!temp_imemload_output_18 & ((\Mux40~15_combout )))))

	.dataa(temp_imemload_output_19),
	.datab(\Mux40~13_combout ),
	.datac(temp_imemload_output_18),
	.datad(\Mux40~15_combout ),
	.cin(gnd),
	.combout(\Mux40~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~16 .lut_mask = 16'hE5E0;
defparam \Mux40~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N9
dffeas \storeregister[8][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][23] .is_wysiwyg = "true";
defparam \storeregister[8][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y39_N3
dffeas \storeregister[10][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][23] .is_wysiwyg = "true";
defparam \storeregister[10][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N2
cycloneive_lcell_comb \Mux40~10 (
// Equation(s):
// \Mux40~10_combout  = (temp_imemload_output_17 & (((\storeregister[10][23]~q ) # (temp_imemload_output_16)))) # (!temp_imemload_output_17 & (\storeregister[8][23]~q  & ((!temp_imemload_output_16))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[8][23]~q ),
	.datac(\storeregister[10][23]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux40~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~10 .lut_mask = 16'hAAE4;
defparam \Mux40~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N20
cycloneive_lcell_comb \Mux40~11 (
// Equation(s):
// \Mux40~11_combout  = (\Mux40~10_combout  & ((\storeregister[11][23]~q ) # ((!temp_imemload_output_16)))) # (!\Mux40~10_combout  & (((\storeregister[9][23]~q  & temp_imemload_output_16))))

	.dataa(\Mux40~10_combout ),
	.datab(\storeregister[11][23]~q ),
	.datac(\storeregister[9][23]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux40~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~11 .lut_mask = 16'hD8AA;
defparam \Mux40~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N12
cycloneive_lcell_comb \Mux41~7 (
// Equation(s):
// \Mux41~7_combout  = (temp_imemload_output_19 & (((\storeregister[27][22]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[19][22]~q  & ((!temp_imemload_output_18))))

	.dataa(\storeregister[19][22]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[27][22]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux41~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~7 .lut_mask = 16'hCCE2;
defparam \Mux41~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N0
cycloneive_lcell_comb \Mux41~8 (
// Equation(s):
// \Mux41~8_combout  = (temp_imemload_output_18 & ((\Mux41~7_combout  & ((\storeregister[31][22]~q ))) # (!\Mux41~7_combout  & (\storeregister[23][22]~q )))) # (!temp_imemload_output_18 & (((\Mux41~7_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[23][22]~q ),
	.datac(\storeregister[31][22]~q ),
	.datad(\Mux41~7_combout ),
	.cin(gnd),
	.combout(\Mux41~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~8 .lut_mask = 16'hF588;
defparam \Mux41~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N15
dffeas \storeregister[20][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][22] .is_wysiwyg = "true";
defparam \storeregister[20][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N14
cycloneive_lcell_comb \Mux41~4 (
// Equation(s):
// \Mux41~4_combout  = (temp_imemload_output_18 & (((\storeregister[20][22]~q ) # (temp_imemload_output_19)))) # (!temp_imemload_output_18 & (\storeregister[16][22]~q  & ((!temp_imemload_output_19))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[16][22]~q ),
	.datac(\storeregister[20][22]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux41~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~4 .lut_mask = 16'hAAE4;
defparam \Mux41~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N18
cycloneive_lcell_comb \Mux41~5 (
// Equation(s):
// \Mux41~5_combout  = (temp_imemload_output_19 & ((\Mux41~4_combout  & ((\storeregister[28][22]~q ))) # (!\Mux41~4_combout  & (\storeregister[24][22]~q )))) # (!temp_imemload_output_19 & (((\Mux41~4_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[24][22]~q ),
	.datac(\storeregister[28][22]~q ),
	.datad(\Mux41~4_combout ),
	.cin(gnd),
	.combout(\Mux41~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~5 .lut_mask = 16'hF588;
defparam \Mux41~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N24
cycloneive_lcell_comb \Mux41~2 (
// Equation(s):
// \Mux41~2_combout  = (temp_imemload_output_18 & (((\storeregister[22][22]~q ) # (temp_imemload_output_19)))) # (!temp_imemload_output_18 & (\storeregister[18][22]~q  & ((!temp_imemload_output_19))))

	.dataa(\storeregister[18][22]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[22][22]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux41~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~2 .lut_mask = 16'hCCE2;
defparam \Mux41~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N30
cycloneive_lcell_comb \Mux41~3 (
// Equation(s):
// \Mux41~3_combout  = (\Mux41~2_combout  & (((\storeregister[30][22]~q ) # (!temp_imemload_output_19)))) # (!\Mux41~2_combout  & (\storeregister[26][22]~q  & ((temp_imemload_output_19))))

	.dataa(\storeregister[26][22]~q ),
	.datab(\Mux41~2_combout ),
	.datac(\storeregister[30][22]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux41~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~3 .lut_mask = 16'hE2CC;
defparam \Mux41~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N30
cycloneive_lcell_comb \Mux41~6 (
// Equation(s):
// \Mux41~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\Mux41~3_combout ))) # (!temp_imemload_output_17 & (\Mux41~5_combout ))))

	.dataa(\Mux41~5_combout ),
	.datab(\Mux41~3_combout ),
	.datac(temp_imemload_output_16),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux41~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~6 .lut_mask = 16'hFC0A;
defparam \Mux41~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N14
cycloneive_lcell_comb \storeregister[21][22]~feeder (
// Equation(s):
// \storeregister[21][22]~feeder_combout  = Mux9

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux9),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[21][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[21][22]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[21][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y34_N15
dffeas \storeregister[21][22] (
	.clk(!CLK),
	.d(\storeregister[21][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[21][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[21][22] .is_wysiwyg = "true";
defparam \storeregister[21][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N26
cycloneive_lcell_comb \Mux41~0 (
// Equation(s):
// \Mux41~0_combout  = (temp_imemload_output_19 & (((\storeregister[25][22]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[17][22]~q  & ((!temp_imemload_output_18))))

	.dataa(\storeregister[17][22]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[25][22]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~0 .lut_mask = 16'hCCE2;
defparam \Mux41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N18
cycloneive_lcell_comb \Mux41~1 (
// Equation(s):
// \Mux41~1_combout  = (\Mux41~0_combout  & ((\storeregister[29][22]~q ) # ((!temp_imemload_output_18)))) # (!\Mux41~0_combout  & (((\storeregister[21][22]~q  & temp_imemload_output_18))))

	.dataa(\storeregister[29][22]~q ),
	.datab(\storeregister[21][22]~q ),
	.datac(\Mux41~0_combout ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~1 .lut_mask = 16'hACF0;
defparam \Mux41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N10
cycloneive_lcell_comb \Mux41~17 (
// Equation(s):
// \Mux41~17_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[13][22]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & (\storeregister[12][22]~q )))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[12][22]~q ),
	.datad(\storeregister[13][22]~q ),
	.cin(gnd),
	.combout(\Mux41~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~17 .lut_mask = 16'hBA98;
defparam \Mux41~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N12
cycloneive_lcell_comb \Mux41~18 (
// Equation(s):
// \Mux41~18_combout  = (\Mux41~17_combout  & (((\storeregister[15][22]~q )) # (!temp_imemload_output_17))) # (!\Mux41~17_combout  & (temp_imemload_output_17 & ((\storeregister[14][22]~q ))))

	.dataa(\Mux41~17_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[15][22]~q ),
	.datad(\storeregister[14][22]~q ),
	.cin(gnd),
	.combout(\Mux41~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~18 .lut_mask = 16'hE6A2;
defparam \Mux41~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N0
cycloneive_lcell_comb \Mux41~10 (
// Equation(s):
// \Mux41~10_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[5][22]~q ))) # (!temp_imemload_output_16 & (\storeregister[4][22]~q ))))

	.dataa(\storeregister[4][22]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][22]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux41~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~10 .lut_mask = 16'hFC22;
defparam \Mux41~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N2
cycloneive_lcell_comb \Mux41~11 (
// Equation(s):
// \Mux41~11_combout  = (\Mux41~10_combout  & (((\storeregister[7][22]~q )) # (!temp_imemload_output_17))) # (!\Mux41~10_combout  & (temp_imemload_output_17 & (\storeregister[6][22]~q )))

	.dataa(\Mux41~10_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[6][22]~q ),
	.datad(\storeregister[7][22]~q ),
	.cin(gnd),
	.combout(\Mux41~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~11 .lut_mask = 16'hEA62;
defparam \Mux41~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y39_N1
dffeas \storeregister[8][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[8][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[8][22] .is_wysiwyg = "true";
defparam \storeregister[8][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N0
cycloneive_lcell_comb \Mux41~12 (
// Equation(s):
// \Mux41~12_combout  = (temp_imemload_output_16 & (temp_imemload_output_17)) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[10][22]~q ))) # (!temp_imemload_output_17 & (\storeregister[8][22]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[8][22]~q ),
	.datad(\storeregister[10][22]~q ),
	.cin(gnd),
	.combout(\Mux41~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~12 .lut_mask = 16'hDC98;
defparam \Mux41~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N22
cycloneive_lcell_comb \Mux41~13 (
// Equation(s):
// \Mux41~13_combout  = (temp_imemload_output_16 & ((\Mux41~12_combout  & ((\storeregister[11][22]~q ))) # (!\Mux41~12_combout  & (\storeregister[9][22]~q )))) # (!temp_imemload_output_16 & (((\Mux41~12_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[9][22]~q ),
	.datac(\storeregister[11][22]~q ),
	.datad(\Mux41~12_combout ),
	.cin(gnd),
	.combout(\Mux41~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~13 .lut_mask = 16'hF588;
defparam \Mux41~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N17
dffeas \storeregister[3][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][22] .is_wysiwyg = "true";
defparam \storeregister[3][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N27
dffeas \storeregister[1][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][22] .is_wysiwyg = "true";
defparam \storeregister[1][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N26
cycloneive_lcell_comb \Mux41~14 (
// Equation(s):
// \Mux41~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][22]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][22]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[3][22]~q ),
	.datac(\storeregister[1][22]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux41~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~14 .lut_mask = 16'hD800;
defparam \Mux41~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N2
cycloneive_lcell_comb \Mux41~15 (
// Equation(s):
// \Mux41~15_combout  = (\Mux41~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][22]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux41~14_combout ),
	.datac(\storeregister[2][22]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux41~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~15 .lut_mask = 16'hCCEC;
defparam \Mux41~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N10
cycloneive_lcell_comb \Mux41~16 (
// Equation(s):
// \Mux41~16_combout  = (temp_imemload_output_19 & ((\Mux41~13_combout ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\Mux41~15_combout  & !temp_imemload_output_18))))

	.dataa(\Mux41~13_combout ),
	.datab(\Mux41~15_combout ),
	.datac(temp_imemload_output_19),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux41~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~16 .lut_mask = 16'hF0AC;
defparam \Mux41~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N0
cycloneive_lcell_comb \Mux42~7 (
// Equation(s):
// \Mux42~7_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[23][21]~q ))) # (!temp_imemload_output_18 & (\storeregister[19][21]~q ))))

	.dataa(\storeregister[19][21]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[23][21]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux42~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~7 .lut_mask = 16'hFC22;
defparam \Mux42~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N6
cycloneive_lcell_comb \Mux42~8 (
// Equation(s):
// \Mux42~8_combout  = (temp_imemload_output_19 & ((\Mux42~7_combout  & (\storeregister[31][21]~q )) # (!\Mux42~7_combout  & ((\storeregister[27][21]~q ))))) # (!temp_imemload_output_19 & (\Mux42~7_combout ))

	.dataa(temp_imemload_output_19),
	.datab(\Mux42~7_combout ),
	.datac(\storeregister[31][21]~q ),
	.datad(\storeregister[27][21]~q ),
	.cin(gnd),
	.combout(\Mux42~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~8 .lut_mask = 16'hE6C4;
defparam \Mux42~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N31
dffeas \storeregister[20][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][21] .is_wysiwyg = "true";
defparam \storeregister[20][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N11
dffeas \storeregister[16][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][21] .is_wysiwyg = "true";
defparam \storeregister[16][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N10
cycloneive_lcell_comb \Mux42~4 (
// Equation(s):
// \Mux42~4_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\storeregister[24][21]~q )) # (!temp_imemload_output_19 & ((\storeregister[16][21]~q )))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[24][21]~q ),
	.datac(\storeregister[16][21]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux42~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~4 .lut_mask = 16'hEE50;
defparam \Mux42~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N4
cycloneive_lcell_comb \Mux42~5 (
// Equation(s):
// \Mux42~5_combout  = (temp_imemload_output_18 & ((\Mux42~4_combout  & (\storeregister[28][21]~q )) # (!\Mux42~4_combout  & ((\storeregister[20][21]~q ))))) # (!temp_imemload_output_18 & (((\Mux42~4_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[28][21]~q ),
	.datac(\storeregister[20][21]~q ),
	.datad(\Mux42~4_combout ),
	.cin(gnd),
	.combout(\Mux42~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~5 .lut_mask = 16'hDDA0;
defparam \Mux42~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N31
dffeas \storeregister[30][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][21] .is_wysiwyg = "true";
defparam \storeregister[30][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N30
cycloneive_lcell_comb \Mux42~3 (
// Equation(s):
// \Mux42~3_combout  = (\Mux42~2_combout  & (((\storeregister[30][21]~q )) # (!temp_imemload_output_18))) # (!\Mux42~2_combout  & (temp_imemload_output_18 & ((\storeregister[22][21]~q ))))

	.dataa(\Mux42~2_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[30][21]~q ),
	.datad(\storeregister[22][21]~q ),
	.cin(gnd),
	.combout(\Mux42~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~3 .lut_mask = 16'hE6A2;
defparam \Mux42~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N20
cycloneive_lcell_comb \Mux42~6 (
// Equation(s):
// \Mux42~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\Mux42~3_combout ))) # (!temp_imemload_output_17 & (\Mux42~5_combout ))))

	.dataa(\Mux42~5_combout ),
	.datab(temp_imemload_output_16),
	.datac(\Mux42~3_combout ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux42~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~6 .lut_mask = 16'hFC22;
defparam \Mux42~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N22
cycloneive_lcell_comb \Mux42~0 (
// Equation(s):
// \Mux42~0_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[21][21]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[17][21]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[21][21]~q ),
	.datad(\storeregister[17][21]~q ),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~0 .lut_mask = 16'hB9A8;
defparam \Mux42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N26
cycloneive_lcell_comb \Mux42~1 (
// Equation(s):
// \Mux42~1_combout  = (temp_imemload_output_19 & ((\Mux42~0_combout  & (\storeregister[29][21]~q )) # (!\Mux42~0_combout  & ((\storeregister[25][21]~q ))))) # (!temp_imemload_output_19 & (((\Mux42~0_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[29][21]~q ),
	.datac(\Mux42~0_combout ),
	.datad(\storeregister[25][21]~q ),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~1 .lut_mask = 16'hDAD0;
defparam \Mux42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N2
cycloneive_lcell_comb \Mux42~14 (
// Equation(s):
// \Mux42~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][21]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][21]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[3][21]~q ),
	.datac(\storeregister[1][21]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux42~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~14 .lut_mask = 16'hD800;
defparam \Mux42~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N31
dffeas \storeregister[2][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[2][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[2][21] .is_wysiwyg = "true";
defparam \storeregister[2][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N30
cycloneive_lcell_comb \Mux42~15 (
// Equation(s):
// \Mux42~15_combout  = (\Mux42~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][21]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux42~14_combout ),
	.datac(\storeregister[2][21]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux42~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~15 .lut_mask = 16'hCCEC;
defparam \Mux42~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N6
cycloneive_lcell_comb \Mux42~12 (
// Equation(s):
// \Mux42~12_combout  = (temp_imemload_output_16 & ((\storeregister[5][21]~q ) # ((temp_imemload_output_17)))) # (!temp_imemload_output_16 & (((\storeregister[4][21]~q  & !temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[5][21]~q ),
	.datac(\storeregister[4][21]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux42~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~12 .lut_mask = 16'hAAD8;
defparam \Mux42~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N4
cycloneive_lcell_comb \Mux42~13 (
// Equation(s):
// \Mux42~13_combout  = (temp_imemload_output_17 & ((\Mux42~12_combout  & (\storeregister[7][21]~q )) # (!\Mux42~12_combout  & ((\storeregister[6][21]~q ))))) # (!temp_imemload_output_17 & (\Mux42~12_combout ))

	.dataa(temp_imemload_output_17),
	.datab(\Mux42~12_combout ),
	.datac(\storeregister[7][21]~q ),
	.datad(\storeregister[6][21]~q ),
	.cin(gnd),
	.combout(\Mux42~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~13 .lut_mask = 16'hE6C4;
defparam \Mux42~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N6
cycloneive_lcell_comb \Mux42~16 (
// Equation(s):
// \Mux42~16_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\Mux42~13_combout ))) # (!temp_imemload_output_18 & (\Mux42~15_combout ))))

	.dataa(\Mux42~15_combout ),
	.datab(temp_imemload_output_19),
	.datac(temp_imemload_output_18),
	.datad(\Mux42~13_combout ),
	.cin(gnd),
	.combout(\Mux42~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~16 .lut_mask = 16'hF2C2;
defparam \Mux42~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N18
cycloneive_lcell_comb \Mux42~17 (
// Equation(s):
// \Mux42~17_combout  = (temp_imemload_output_16 & ((\storeregister[13][21]~q ) # ((temp_imemload_output_17)))) # (!temp_imemload_output_16 & (((\storeregister[12][21]~q  & !temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[13][21]~q ),
	.datac(\storeregister[12][21]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux42~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~17 .lut_mask = 16'hAAD8;
defparam \Mux42~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N0
cycloneive_lcell_comb \Mux42~18 (
// Equation(s):
// \Mux42~18_combout  = (temp_imemload_output_17 & ((\Mux42~17_combout  & (\storeregister[15][21]~q )) # (!\Mux42~17_combout  & ((\storeregister[14][21]~q ))))) # (!temp_imemload_output_17 & (((\Mux42~17_combout ))))

	.dataa(\storeregister[15][21]~q ),
	.datab(temp_imemload_output_17),
	.datac(\Mux42~17_combout ),
	.datad(\storeregister[14][21]~q ),
	.cin(gnd),
	.combout(\Mux42~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~18 .lut_mask = 16'hBCB0;
defparam \Mux42~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y39_N13
dffeas \storeregister[9][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[9][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[9][21] .is_wysiwyg = "true";
defparam \storeregister[9][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N0
cycloneive_lcell_comb \Mux42~10 (
// Equation(s):
// \Mux42~10_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[10][21]~q ))) # (!temp_imemload_output_17 & (\storeregister[8][21]~q ))))

	.dataa(\storeregister[8][21]~q ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[10][21]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux42~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~10 .lut_mask = 16'hFC22;
defparam \Mux42~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N12
cycloneive_lcell_comb \Mux42~11 (
// Equation(s):
// \Mux42~11_combout  = (temp_imemload_output_16 & ((\Mux42~10_combout  & (\storeregister[11][21]~q )) # (!\Mux42~10_combout  & ((\storeregister[9][21]~q ))))) # (!temp_imemload_output_16 & (((\Mux42~10_combout ))))

	.dataa(\storeregister[11][21]~q ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[9][21]~q ),
	.datad(\Mux42~10_combout ),
	.cin(gnd),
	.combout(\Mux42~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~11 .lut_mask = 16'hBBC0;
defparam \Mux42~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N4
cycloneive_lcell_comb \Mux43~0 (
// Equation(s):
// \Mux43~0_combout  = (temp_imemload_output_19 & (((\storeregister[25][20]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[17][20]~q  & ((!temp_imemload_output_18))))

	.dataa(\storeregister[17][20]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[25][20]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~0 .lut_mask = 16'hCCE2;
defparam \Mux43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N6
cycloneive_lcell_comb \Mux43~1 (
// Equation(s):
// \Mux43~1_combout  = (temp_imemload_output_18 & ((\Mux43~0_combout  & ((\storeregister[29][20]~q ))) # (!\Mux43~0_combout  & (\storeregister[21][20]~q )))) # (!temp_imemload_output_18 & (\Mux43~0_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux43~0_combout ),
	.datac(\storeregister[21][20]~q ),
	.datad(\storeregister[29][20]~q ),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~1 .lut_mask = 16'hEC64;
defparam \Mux43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N20
cycloneive_lcell_comb \Mux43~3 (
// Equation(s):
// \Mux43~3_combout  = (\Mux43~2_combout  & (((\storeregister[30][20]~q ) # (!temp_imemload_output_19)))) # (!\Mux43~2_combout  & (\storeregister[26][20]~q  & ((temp_imemload_output_19))))

	.dataa(\Mux43~2_combout ),
	.datab(\storeregister[26][20]~q ),
	.datac(\storeregister[30][20]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux43~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~3 .lut_mask = 16'hE4AA;
defparam \Mux43~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N4
cycloneive_lcell_comb \Mux43~4 (
// Equation(s):
// \Mux43~4_combout  = (temp_imemload_output_18 & (((\storeregister[20][20]~q ) # (temp_imemload_output_19)))) # (!temp_imemload_output_18 & (\storeregister[16][20]~q  & ((!temp_imemload_output_19))))

	.dataa(\storeregister[16][20]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[20][20]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux43~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~4 .lut_mask = 16'hCCE2;
defparam \Mux43~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N3
dffeas \storeregister[24][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][20] .is_wysiwyg = "true";
defparam \storeregister[24][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N2
cycloneive_lcell_comb \Mux43~5 (
// Equation(s):
// \Mux43~5_combout  = (temp_imemload_output_19 & ((\Mux43~4_combout  & ((\storeregister[28][20]~q ))) # (!\Mux43~4_combout  & (\storeregister[24][20]~q )))) # (!temp_imemload_output_19 & (\Mux43~4_combout ))

	.dataa(temp_imemload_output_19),
	.datab(\Mux43~4_combout ),
	.datac(\storeregister[24][20]~q ),
	.datad(\storeregister[28][20]~q ),
	.cin(gnd),
	.combout(\Mux43~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~5 .lut_mask = 16'hEC64;
defparam \Mux43~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N30
cycloneive_lcell_comb \Mux43~6 (
// Equation(s):
// \Mux43~6_combout  = (temp_imemload_output_17 & ((\Mux43~3_combout ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((\Mux43~5_combout  & !temp_imemload_output_16))))

	.dataa(temp_imemload_output_17),
	.datab(\Mux43~3_combout ),
	.datac(\Mux43~5_combout ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux43~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~6 .lut_mask = 16'hAAD8;
defparam \Mux43~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N8
cycloneive_lcell_comb \storeregister[23][20]~feeder (
// Equation(s):
// \storeregister[23][20]~feeder_combout  = Mux11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux11),
	.cin(gnd),
	.combout(\storeregister[23][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[23][20]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[23][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N9
dffeas \storeregister[23][20] (
	.clk(!CLK),
	.d(\storeregister[23][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[23][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[23][20] .is_wysiwyg = "true";
defparam \storeregister[23][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N20
cycloneive_lcell_comb \Mux43~7 (
// Equation(s):
// \Mux43~7_combout  = (temp_imemload_output_19 & (((\storeregister[27][20]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[19][20]~q  & ((!temp_imemload_output_18))))

	.dataa(\storeregister[19][20]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[27][20]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux43~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~7 .lut_mask = 16'hCCE2;
defparam \Mux43~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N10
cycloneive_lcell_comb \Mux43~8 (
// Equation(s):
// \Mux43~8_combout  = (temp_imemload_output_18 & ((\Mux43~7_combout  & ((\storeregister[31][20]~q ))) # (!\Mux43~7_combout  & (\storeregister[23][20]~q )))) # (!temp_imemload_output_18 & (((\Mux43~7_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[23][20]~q ),
	.datac(\storeregister[31][20]~q ),
	.datad(\Mux43~7_combout ),
	.cin(gnd),
	.combout(\Mux43~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~8 .lut_mask = 16'hF588;
defparam \Mux43~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N8
cycloneive_lcell_comb \Mux43~10 (
// Equation(s):
// \Mux43~10_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][20]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & ((\storeregister[4][20]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][20]~q ),
	.datad(\storeregister[4][20]~q ),
	.cin(gnd),
	.combout(\Mux43~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~10 .lut_mask = 16'hB9A8;
defparam \Mux43~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N8
cycloneive_lcell_comb \Mux43~11 (
// Equation(s):
// \Mux43~11_combout  = (temp_imemload_output_17 & ((\Mux43~10_combout  & (\storeregister[7][20]~q )) # (!\Mux43~10_combout  & ((\storeregister[6][20]~q ))))) # (!temp_imemload_output_17 & (((\Mux43~10_combout ))))

	.dataa(\storeregister[7][20]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[6][20]~q ),
	.datad(\Mux43~10_combout ),
	.cin(gnd),
	.combout(\Mux43~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~11 .lut_mask = 16'hBBC0;
defparam \Mux43~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y41_N31
dffeas \storeregister[1][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][20] .is_wysiwyg = "true";
defparam \storeregister[1][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N29
dffeas \storeregister[3][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][20] .is_wysiwyg = "true";
defparam \storeregister[3][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N30
cycloneive_lcell_comb \Mux43~14 (
// Equation(s):
// \Mux43~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[3][20]~q ))) # (!temp_imemload_output_17 & (\storeregister[1][20]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[1][20]~q ),
	.datad(\storeregister[3][20]~q ),
	.cin(gnd),
	.combout(\Mux43~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~14 .lut_mask = 16'hA820;
defparam \Mux43~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N28
cycloneive_lcell_comb \Mux43~15 (
// Equation(s):
// \Mux43~15_combout  = (\Mux43~14_combout ) # ((!temp_imemload_output_16 & (temp_imemload_output_17 & \storeregister[2][20]~q )))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[2][20]~q ),
	.datad(\Mux43~14_combout ),
	.cin(gnd),
	.combout(\Mux43~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~15 .lut_mask = 16'hFF40;
defparam \Mux43~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N8
cycloneive_lcell_comb \Mux43~12 (
// Equation(s):
// \Mux43~12_combout  = (temp_imemload_output_17 & ((\storeregister[10][20]~q ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((\storeregister[8][20]~q  & !temp_imemload_output_16))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[10][20]~q ),
	.datac(\storeregister[8][20]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux43~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~12 .lut_mask = 16'hAAD8;
defparam \Mux43~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N18
cycloneive_lcell_comb \Mux43~13 (
// Equation(s):
// \Mux43~13_combout  = (temp_imemload_output_16 & ((\Mux43~12_combout  & ((\storeregister[11][20]~q ))) # (!\Mux43~12_combout  & (\storeregister[9][20]~q )))) # (!temp_imemload_output_16 & (((\Mux43~12_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[9][20]~q ),
	.datac(\storeregister[11][20]~q ),
	.datad(\Mux43~12_combout ),
	.cin(gnd),
	.combout(\Mux43~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~13 .lut_mask = 16'hF588;
defparam \Mux43~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N2
cycloneive_lcell_comb \Mux43~16 (
// Equation(s):
// \Mux43~16_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\Mux43~13_combout ))) # (!temp_imemload_output_19 & (\Mux43~15_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\Mux43~15_combout ),
	.datac(temp_imemload_output_19),
	.datad(\Mux43~13_combout ),
	.cin(gnd),
	.combout(\Mux43~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~16 .lut_mask = 16'hF4A4;
defparam \Mux43~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N20
cycloneive_lcell_comb \Mux43~17 (
// Equation(s):
// \Mux43~17_combout  = (temp_imemload_output_16 & (((\storeregister[13][20]~q ) # (temp_imemload_output_17)))) # (!temp_imemload_output_16 & (\storeregister[12][20]~q  & ((!temp_imemload_output_17))))

	.dataa(\storeregister[12][20]~q ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[13][20]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux43~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~17 .lut_mask = 16'hCCE2;
defparam \Mux43~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N24
cycloneive_lcell_comb \Mux43~18 (
// Equation(s):
// \Mux43~18_combout  = (temp_imemload_output_17 & ((\Mux43~17_combout  & (\storeregister[15][20]~q )) # (!\Mux43~17_combout  & ((\storeregister[14][20]~q ))))) # (!temp_imemload_output_17 & (((\Mux43~17_combout ))))

	.dataa(\storeregister[15][20]~q ),
	.datab(temp_imemload_output_17),
	.datac(\Mux43~17_combout ),
	.datad(\storeregister[14][20]~q ),
	.cin(gnd),
	.combout(\Mux43~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~18 .lut_mask = 16'hBCB0;
defparam \Mux43~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N6
cycloneive_lcell_comb \Mux44~7 (
// Equation(s):
// \Mux44~7_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\storeregister[23][19]~q )) # (!temp_imemload_output_18 & ((\storeregister[19][19]~q )))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[23][19]~q ),
	.datad(\storeregister[19][19]~q ),
	.cin(gnd),
	.combout(\Mux44~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~7 .lut_mask = 16'hD9C8;
defparam \Mux44~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N24
cycloneive_lcell_comb \Mux44~8 (
// Equation(s):
// \Mux44~8_combout  = (temp_imemload_output_19 & ((\Mux44~7_combout  & ((\storeregister[31][19]~q ))) # (!\Mux44~7_combout  & (\storeregister[27][19]~q )))) # (!temp_imemload_output_19 & (((\Mux44~7_combout ))))

	.dataa(\storeregister[27][19]~q ),
	.datab(\storeregister[31][19]~q ),
	.datac(temp_imemload_output_19),
	.datad(\Mux44~7_combout ),
	.cin(gnd),
	.combout(\Mux44~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~8 .lut_mask = 16'hCFA0;
defparam \Mux44~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N30
cycloneive_lcell_comb \Mux44~0 (
// Equation(s):
// \Mux44~0_combout  = (temp_imemload_output_18 & ((\storeregister[21][19]~q ) # ((temp_imemload_output_19)))) # (!temp_imemload_output_18 & (((\storeregister[17][19]~q  & !temp_imemload_output_19))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[21][19]~q ),
	.datac(\storeregister[17][19]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~0 .lut_mask = 16'hAAD8;
defparam \Mux44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N10
cycloneive_lcell_comb \Mux44~1 (
// Equation(s):
// \Mux44~1_combout  = (temp_imemload_output_19 & ((\Mux44~0_combout  & (\storeregister[29][19]~q )) # (!\Mux44~0_combout  & ((\storeregister[25][19]~q ))))) # (!temp_imemload_output_19 & (\Mux44~0_combout ))

	.dataa(temp_imemload_output_19),
	.datab(\Mux44~0_combout ),
	.datac(\storeregister[29][19]~q ),
	.datad(\storeregister[25][19]~q ),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~1 .lut_mask = 16'hE6C4;
defparam \Mux44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N4
cycloneive_lcell_comb \storeregister[26][19]~feeder (
// Equation(s):
// \storeregister[26][19]~feeder_combout  = Mux12

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux12),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[26][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[26][19]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[26][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N5
dffeas \storeregister[26][19] (
	.clk(!CLK),
	.d(\storeregister[26][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[26][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[26][19] .is_wysiwyg = "true";
defparam \storeregister[26][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N6
cycloneive_lcell_comb \Mux44~2 (
// Equation(s):
// \Mux44~2_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[26][19]~q ))) # (!temp_imemload_output_19 & (\storeregister[18][19]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[18][19]~q ),
	.datad(\storeregister[26][19]~q ),
	.cin(gnd),
	.combout(\Mux44~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~2 .lut_mask = 16'hDC98;
defparam \Mux44~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N8
cycloneive_lcell_comb \Mux44~3 (
// Equation(s):
// \Mux44~3_combout  = (temp_imemload_output_18 & ((\Mux44~2_combout  & (\storeregister[30][19]~q )) # (!\Mux44~2_combout  & ((\storeregister[22][19]~q ))))) # (!temp_imemload_output_18 & (((\Mux44~2_combout ))))

	.dataa(\storeregister[30][19]~q ),
	.datab(temp_imemload_output_18),
	.datac(\Mux44~2_combout ),
	.datad(\storeregister[22][19]~q ),
	.cin(gnd),
	.combout(\Mux44~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~3 .lut_mask = 16'hBCB0;
defparam \Mux44~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N20
cycloneive_lcell_comb \storeregister[24][19]~feeder (
// Equation(s):
// \storeregister[24][19]~feeder_combout  = Mux12

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux12),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[24][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][19]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[24][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N21
dffeas \storeregister[24][19] (
	.clk(!CLK),
	.d(\storeregister[24][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][19] .is_wysiwyg = "true";
defparam \storeregister[24][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N10
cycloneive_lcell_comb \Mux44~4 (
// Equation(s):
// \Mux44~4_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\storeregister[24][19]~q )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & (\storeregister[16][19]~q )))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[16][19]~q ),
	.datad(\storeregister[24][19]~q ),
	.cin(gnd),
	.combout(\Mux44~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~4 .lut_mask = 16'hBA98;
defparam \Mux44~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N18
cycloneive_lcell_comb \Mux44~5 (
// Equation(s):
// \Mux44~5_combout  = (temp_imemload_output_18 & ((\Mux44~4_combout  & (\storeregister[28][19]~q )) # (!\Mux44~4_combout  & ((\storeregister[20][19]~q ))))) # (!temp_imemload_output_18 & (((\Mux44~4_combout ))))

	.dataa(\storeregister[28][19]~q ),
	.datab(temp_imemload_output_18),
	.datac(\Mux44~4_combout ),
	.datad(\storeregister[20][19]~q ),
	.cin(gnd),
	.combout(\Mux44~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~5 .lut_mask = 16'hBCB0;
defparam \Mux44~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N12
cycloneive_lcell_comb \Mux44~6 (
// Equation(s):
// \Mux44~6_combout  = (temp_imemload_output_16 & (temp_imemload_output_17)) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\Mux44~3_combout )) # (!temp_imemload_output_17 & ((\Mux44~5_combout )))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\Mux44~3_combout ),
	.datad(\Mux44~5_combout ),
	.cin(gnd),
	.combout(\Mux44~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~6 .lut_mask = 16'hD9C8;
defparam \Mux44~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y39_N29
dffeas \storeregister[10][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][19] .is_wysiwyg = "true";
defparam \storeregister[10][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N28
cycloneive_lcell_comb \Mux44~10 (
// Equation(s):
// \Mux44~10_combout  = (temp_imemload_output_17 & (((\storeregister[10][19]~q ) # (temp_imemload_output_16)))) # (!temp_imemload_output_17 & (\storeregister[8][19]~q  & ((!temp_imemload_output_16))))

	.dataa(\storeregister[8][19]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[10][19]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux44~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~10 .lut_mask = 16'hCCE2;
defparam \Mux44~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N24
cycloneive_lcell_comb \Mux44~11 (
// Equation(s):
// \Mux44~11_combout  = (temp_imemload_output_16 & ((\Mux44~10_combout  & ((\storeregister[11][19]~q ))) # (!\Mux44~10_combout  & (\storeregister[9][19]~q )))) # (!temp_imemload_output_16 & (\Mux44~10_combout ))

	.dataa(temp_imemload_output_16),
	.datab(\Mux44~10_combout ),
	.datac(\storeregister[9][19]~q ),
	.datad(\storeregister[11][19]~q ),
	.cin(gnd),
	.combout(\Mux44~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~11 .lut_mask = 16'hEC64;
defparam \Mux44~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N18
cycloneive_lcell_comb \Mux44~14 (
// Equation(s):
// \Mux44~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][19]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][19]~q )))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[3][19]~q ),
	.datac(\storeregister[1][19]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux44~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~14 .lut_mask = 16'h88A0;
defparam \Mux44~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N14
cycloneive_lcell_comb \Mux44~15 (
// Equation(s):
// \Mux44~15_combout  = (\Mux44~14_combout ) # ((!temp_imemload_output_16 & (\storeregister[2][19]~q  & temp_imemload_output_17)))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[2][19]~q ),
	.datac(temp_imemload_output_17),
	.datad(\Mux44~14_combout ),
	.cin(gnd),
	.combout(\Mux44~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~15 .lut_mask = 16'hFF40;
defparam \Mux44~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y40_N23
dffeas \storeregister[4][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][19] .is_wysiwyg = "true";
defparam \storeregister[4][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y40_N22
cycloneive_lcell_comb \Mux44~12 (
// Equation(s):
// \Mux44~12_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][19]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & (\storeregister[4][19]~q )))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[4][19]~q ),
	.datad(\storeregister[5][19]~q ),
	.cin(gnd),
	.combout(\Mux44~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~12 .lut_mask = 16'hBA98;
defparam \Mux44~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N26
cycloneive_lcell_comb \Mux44~13 (
// Equation(s):
// \Mux44~13_combout  = (temp_imemload_output_17 & ((\Mux44~12_combout  & ((\storeregister[7][19]~q ))) # (!\Mux44~12_combout  & (\storeregister[6][19]~q )))) # (!temp_imemload_output_17 & (((\Mux44~12_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[6][19]~q ),
	.datac(\storeregister[7][19]~q ),
	.datad(\Mux44~12_combout ),
	.cin(gnd),
	.combout(\Mux44~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~13 .lut_mask = 16'hF588;
defparam \Mux44~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N4
cycloneive_lcell_comb \Mux44~16 (
// Equation(s):
// \Mux44~16_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19) # (\Mux44~13_combout )))) # (!temp_imemload_output_18 & (\Mux44~15_combout  & (!temp_imemload_output_19)))

	.dataa(\Mux44~15_combout ),
	.datab(temp_imemload_output_18),
	.datac(temp_imemload_output_19),
	.datad(\Mux44~13_combout ),
	.cin(gnd),
	.combout(\Mux44~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~16 .lut_mask = 16'hCEC2;
defparam \Mux44~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N4
cycloneive_lcell_comb \Mux44~17 (
// Equation(s):
// \Mux44~17_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][19]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][19]~q ))))

	.dataa(\storeregister[12][19]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[13][19]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux44~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~17 .lut_mask = 16'hFC22;
defparam \Mux44~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N16
cycloneive_lcell_comb \Mux44~18 (
// Equation(s):
// \Mux44~18_combout  = (\Mux44~17_combout  & ((\storeregister[15][19]~q ) # ((!temp_imemload_output_17)))) # (!\Mux44~17_combout  & (((\storeregister[14][19]~q  & temp_imemload_output_17))))

	.dataa(\Mux44~17_combout ),
	.datab(\storeregister[15][19]~q ),
	.datac(\storeregister[14][19]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux44~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~18 .lut_mask = 16'hD8AA;
defparam \Mux44~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N23
dffeas \storeregister[18][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[18][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[18][10] .is_wysiwyg = "true";
defparam \storeregister[18][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N22
cycloneive_lcell_comb \Mux53~2 (
// Equation(s):
// \Mux53~2_combout  = (temp_imemload_output_19 & ((\storeregister[26][10]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\storeregister[18][10]~q  & !temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[26][10]~q ),
	.datac(\storeregister[18][10]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux53~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~2 .lut_mask = 16'hAAD8;
defparam \Mux53~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N0
cycloneive_lcell_comb \Mux53~3 (
// Equation(s):
// \Mux53~3_combout  = (temp_imemload_output_18 & ((\Mux53~2_combout  & ((\storeregister[30][10]~q ))) # (!\Mux53~2_combout  & (\storeregister[22][10]~q )))) # (!temp_imemload_output_18 & (((\Mux53~2_combout ))))

	.dataa(\storeregister[22][10]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[30][10]~q ),
	.datad(\Mux53~2_combout ),
	.cin(gnd),
	.combout(\Mux53~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~3 .lut_mask = 16'hF388;
defparam \Mux53~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N1
dffeas \storeregister[16][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][10] .is_wysiwyg = "true";
defparam \storeregister[16][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N31
dffeas \storeregister[24][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][10] .is_wysiwyg = "true";
defparam \storeregister[24][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N30
cycloneive_lcell_comb \Mux53~4 (
// Equation(s):
// \Mux53~4_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[24][10]~q ))) # (!temp_imemload_output_19 & (\storeregister[16][10]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[16][10]~q ),
	.datac(\storeregister[24][10]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux53~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~4 .lut_mask = 16'hFA44;
defparam \Mux53~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N24
cycloneive_lcell_comb \Mux53~5 (
// Equation(s):
// \Mux53~5_combout  = (temp_imemload_output_18 & ((\Mux53~4_combout  & ((\storeregister[28][10]~q ))) # (!\Mux53~4_combout  & (\storeregister[20][10]~q )))) # (!temp_imemload_output_18 & (\Mux53~4_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux53~4_combout ),
	.datac(\storeregister[20][10]~q ),
	.datad(\storeregister[28][10]~q ),
	.cin(gnd),
	.combout(\Mux53~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~5 .lut_mask = 16'hEC64;
defparam \Mux53~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N26
cycloneive_lcell_comb \Mux53~6 (
// Equation(s):
// \Mux53~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\Mux53~3_combout )) # (!temp_imemload_output_17 & ((\Mux53~5_combout )))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux53~3_combout ),
	.datac(\Mux53~5_combout ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux53~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~6 .lut_mask = 16'hEE50;
defparam \Mux53~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N12
cycloneive_lcell_comb \Mux53~7 (
// Equation(s):
// \Mux53~7_combout  = (temp_imemload_output_18 & (((\storeregister[23][10]~q ) # (temp_imemload_output_19)))) # (!temp_imemload_output_18 & (\storeregister[19][10]~q  & ((!temp_imemload_output_19))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[19][10]~q ),
	.datac(\storeregister[23][10]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux53~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~7 .lut_mask = 16'hAAE4;
defparam \Mux53~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N24
cycloneive_lcell_comb \Mux53~8 (
// Equation(s):
// \Mux53~8_combout  = (\Mux53~7_combout  & ((\storeregister[31][10]~q ) # ((!temp_imemload_output_19)))) # (!\Mux53~7_combout  & (((temp_imemload_output_19 & \storeregister[27][10]~q ))))

	.dataa(\Mux53~7_combout ),
	.datab(\storeregister[31][10]~q ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[27][10]~q ),
	.cin(gnd),
	.combout(\Mux53~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~8 .lut_mask = 16'hDA8A;
defparam \Mux53~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N8
cycloneive_lcell_comb \Mux53~0 (
// Equation(s):
// \Mux53~0_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[21][10]~q ))) # (!temp_imemload_output_18 & (\storeregister[17][10]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[17][10]~q ),
	.datad(\storeregister[21][10]~q ),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~0 .lut_mask = 16'hDC98;
defparam \Mux53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N24
cycloneive_lcell_comb \Mux53~1 (
// Equation(s):
// \Mux53~1_combout  = (temp_imemload_output_19 & ((\Mux53~0_combout  & (\storeregister[29][10]~q )) # (!\Mux53~0_combout  & ((\storeregister[25][10]~q ))))) # (!temp_imemload_output_19 & (\Mux53~0_combout ))

	.dataa(temp_imemload_output_19),
	.datab(\Mux53~0_combout ),
	.datac(\storeregister[29][10]~q ),
	.datad(\storeregister[25][10]~q ),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~1 .lut_mask = 16'hE6C4;
defparam \Mux53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N12
cycloneive_lcell_comb \Mux53~17 (
// Equation(s):
// \Mux53~17_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][10]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][10]~q ))))

	.dataa(\storeregister[12][10]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[13][10]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux53~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~17 .lut_mask = 16'hFC22;
defparam \Mux53~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N30
cycloneive_lcell_comb \Mux53~18 (
// Equation(s):
// \Mux53~18_combout  = (\Mux53~17_combout  & (((\storeregister[15][10]~q ) # (!temp_imemload_output_17)))) # (!\Mux53~17_combout  & (\storeregister[14][10]~q  & ((temp_imemload_output_17))))

	.dataa(\Mux53~17_combout ),
	.datab(\storeregister[14][10]~q ),
	.datac(\storeregister[15][10]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux53~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~18 .lut_mask = 16'hE4AA;
defparam \Mux53~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N24
cycloneive_lcell_comb \Mux53~10 (
// Equation(s):
// \Mux53~10_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[10][10]~q ))) # (!temp_imemload_output_17 & (\storeregister[8][10]~q ))))

	.dataa(\storeregister[8][10]~q ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[10][10]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux53~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~10 .lut_mask = 16'hFC22;
defparam \Mux53~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N0
cycloneive_lcell_comb \Mux53~11 (
// Equation(s):
// \Mux53~11_combout  = (\Mux53~10_combout  & (((\storeregister[11][10]~q ) # (!temp_imemload_output_16)))) # (!\Mux53~10_combout  & (\storeregister[9][10]~q  & ((temp_imemload_output_16))))

	.dataa(\Mux53~10_combout ),
	.datab(\storeregister[9][10]~q ),
	.datac(\storeregister[11][10]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux53~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~11 .lut_mask = 16'hE4AA;
defparam \Mux53~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y39_N13
dffeas \storeregister[6][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[6][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[6][10] .is_wysiwyg = "true";
defparam \storeregister[6][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y41_N18
cycloneive_lcell_comb \Mux53~12 (
// Equation(s):
// \Mux53~12_combout  = (temp_imemload_output_16 & ((\storeregister[5][10]~q ) # ((temp_imemload_output_17)))) # (!temp_imemload_output_16 & (((\storeregister[4][10]~q  & !temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[5][10]~q ),
	.datac(\storeregister[4][10]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux53~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~12 .lut_mask = 16'hAAD8;
defparam \Mux53~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N12
cycloneive_lcell_comb \Mux53~13 (
// Equation(s):
// \Mux53~13_combout  = (temp_imemload_output_17 & ((\Mux53~12_combout  & (\storeregister[7][10]~q )) # (!\Mux53~12_combout  & ((\storeregister[6][10]~q ))))) # (!temp_imemload_output_17 & (((\Mux53~12_combout ))))

	.dataa(\storeregister[7][10]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[6][10]~q ),
	.datad(\Mux53~12_combout ),
	.cin(gnd),
	.combout(\Mux53~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~13 .lut_mask = 16'hBBC0;
defparam \Mux53~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N31
dffeas \storeregister[1][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][10] .is_wysiwyg = "true";
defparam \storeregister[1][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N30
cycloneive_lcell_comb \Mux53~14 (
// Equation(s):
// \Mux53~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][10]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][10]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[3][10]~q ),
	.datac(\storeregister[1][10]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux53~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~14 .lut_mask = 16'hD800;
defparam \Mux53~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N28
cycloneive_lcell_comb \Mux53~15 (
// Equation(s):
// \Mux53~15_combout  = (\Mux53~14_combout ) # ((!temp_imemload_output_16 & (\storeregister[2][10]~q  & temp_imemload_output_17)))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[2][10]~q ),
	.datac(\Mux53~14_combout ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux53~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~15 .lut_mask = 16'hF4F0;
defparam \Mux53~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N18
cycloneive_lcell_comb \Mux53~16 (
// Equation(s):
// \Mux53~16_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\Mux53~13_combout )) # (!temp_imemload_output_18 & ((\Mux53~15_combout )))))

	.dataa(\Mux53~13_combout ),
	.datab(\Mux53~15_combout ),
	.datac(temp_imemload_output_19),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux53~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~16 .lut_mask = 16'hFA0C;
defparam \Mux53~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N26
cycloneive_lcell_comb \Mux49~7 (
// Equation(s):
// \Mux49~7_combout  = (temp_imemload_output_19 & ((\storeregister[27][14]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\storeregister[19][14]~q  & !temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[27][14]~q ),
	.datac(\storeregister[19][14]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux49~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~7 .lut_mask = 16'hAAD8;
defparam \Mux49~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N28
cycloneive_lcell_comb \Mux49~8 (
// Equation(s):
// \Mux49~8_combout  = (temp_imemload_output_18 & ((\Mux49~7_combout  & ((\storeregister[31][14]~q ))) # (!\Mux49~7_combout  & (\storeregister[23][14]~q )))) # (!temp_imemload_output_18 & (((\Mux49~7_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[23][14]~q ),
	.datac(\Mux49~7_combout ),
	.datad(\storeregister[31][14]~q ),
	.cin(gnd),
	.combout(\Mux49~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~8 .lut_mask = 16'hF858;
defparam \Mux49~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N2
cycloneive_lcell_comb \Mux49~0 (
// Equation(s):
// \Mux49~0_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\storeregister[25][14]~q )) # (!temp_imemload_output_19 & ((\storeregister[17][14]~q )))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[25][14]~q ),
	.datad(\storeregister[17][14]~q ),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~0 .lut_mask = 16'hD9C8;
defparam \Mux49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N30
cycloneive_lcell_comb \Mux49~1 (
// Equation(s):
// \Mux49~1_combout  = (\Mux49~0_combout  & (((\storeregister[29][14]~q )) # (!temp_imemload_output_18))) # (!\Mux49~0_combout  & (temp_imemload_output_18 & ((\storeregister[21][14]~q ))))

	.dataa(\Mux49~0_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[29][14]~q ),
	.datad(\storeregister[21][14]~q ),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~1 .lut_mask = 16'hE6A2;
defparam \Mux49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N18
cycloneive_lcell_comb \Mux49~2 (
// Equation(s):
// \Mux49~2_combout  = (temp_imemload_output_18 & (((\storeregister[22][14]~q ) # (temp_imemload_output_19)))) # (!temp_imemload_output_18 & (\storeregister[18][14]~q  & ((!temp_imemload_output_19))))

	.dataa(\storeregister[18][14]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[22][14]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux49~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~2 .lut_mask = 16'hCCE2;
defparam \Mux49~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N4
cycloneive_lcell_comb \Mux49~3 (
// Equation(s):
// \Mux49~3_combout  = (temp_imemload_output_19 & ((\Mux49~2_combout  & ((\storeregister[30][14]~q ))) # (!\Mux49~2_combout  & (\storeregister[26][14]~q )))) # (!temp_imemload_output_19 & (((\Mux49~2_combout ))))

	.dataa(\storeregister[26][14]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[30][14]~q ),
	.datad(\Mux49~2_combout ),
	.cin(gnd),
	.combout(\Mux49~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~3 .lut_mask = 16'hF388;
defparam \Mux49~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N12
cycloneive_lcell_comb \Mux49~5 (
// Equation(s):
// \Mux49~5_combout  = (\Mux49~4_combout  & (((\storeregister[28][14]~q )) # (!temp_imemload_output_19))) # (!\Mux49~4_combout  & (temp_imemload_output_19 & ((\storeregister[24][14]~q ))))

	.dataa(\Mux49~4_combout ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[28][14]~q ),
	.datad(\storeregister[24][14]~q ),
	.cin(gnd),
	.combout(\Mux49~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~5 .lut_mask = 16'hE6A2;
defparam \Mux49~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N22
cycloneive_lcell_comb \Mux49~6 (
// Equation(s):
// \Mux49~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\Mux49~3_combout )) # (!temp_imemload_output_17 & ((\Mux49~5_combout )))))

	.dataa(\Mux49~3_combout ),
	.datab(temp_imemload_output_16),
	.datac(\Mux49~5_combout ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux49~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~6 .lut_mask = 16'hEE30;
defparam \Mux49~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N18
cycloneive_lcell_comb \Mux49~17 (
// Equation(s):
// \Mux49~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][14]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][14]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[12][14]~q ),
	.datad(\storeregister[13][14]~q ),
	.cin(gnd),
	.combout(\Mux49~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~17 .lut_mask = 16'hDC98;
defparam \Mux49~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N14
cycloneive_lcell_comb \Mux49~18 (
// Equation(s):
// \Mux49~18_combout  = (\Mux49~17_combout  & (((\storeregister[15][14]~q ) # (!temp_imemload_output_17)))) # (!\Mux49~17_combout  & (\storeregister[14][14]~q  & ((temp_imemload_output_17))))

	.dataa(\Mux49~17_combout ),
	.datab(\storeregister[14][14]~q ),
	.datac(\storeregister[15][14]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux49~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~18 .lut_mask = 16'hE4AA;
defparam \Mux49~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N22
cycloneive_lcell_comb \Mux49~12 (
// Equation(s):
// \Mux49~12_combout  = (temp_imemload_output_17 & ((\storeregister[10][14]~q ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((!temp_imemload_output_16 & \storeregister[8][14]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[10][14]~q ),
	.datac(temp_imemload_output_16),
	.datad(\storeregister[8][14]~q ),
	.cin(gnd),
	.combout(\Mux49~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~12 .lut_mask = 16'hADA8;
defparam \Mux49~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N16
cycloneive_lcell_comb \Mux49~13 (
// Equation(s):
// \Mux49~13_combout  = (temp_imemload_output_16 & ((\Mux49~12_combout  & ((\storeregister[11][14]~q ))) # (!\Mux49~12_combout  & (\storeregister[9][14]~q )))) # (!temp_imemload_output_16 & (((\Mux49~12_combout ))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[9][14]~q ),
	.datac(\storeregister[11][14]~q ),
	.datad(\Mux49~12_combout ),
	.cin(gnd),
	.combout(\Mux49~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~13 .lut_mask = 16'hF588;
defparam \Mux49~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N9
dffeas \storeregister[3][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][14] .is_wysiwyg = "true";
defparam \storeregister[3][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N7
dffeas \storeregister[1][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][14] .is_wysiwyg = "true";
defparam \storeregister[1][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N8
cycloneive_lcell_comb \Mux49~14 (
// Equation(s):
// \Mux49~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][14]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][14]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[3][14]~q ),
	.datad(\storeregister[1][14]~q ),
	.cin(gnd),
	.combout(\Mux49~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~14 .lut_mask = 16'hC480;
defparam \Mux49~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N14
cycloneive_lcell_comb \Mux49~15 (
// Equation(s):
// \Mux49~15_combout  = (\Mux49~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][14]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux49~14_combout ),
	.datac(\storeregister[2][14]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux49~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~15 .lut_mask = 16'hCCEC;
defparam \Mux49~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N26
cycloneive_lcell_comb \Mux49~16 (
// Equation(s):
// \Mux49~16_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\Mux49~13_combout )) # (!temp_imemload_output_19 & ((\Mux49~15_combout )))))

	.dataa(\Mux49~13_combout ),
	.datab(temp_imemload_output_18),
	.datac(temp_imemload_output_19),
	.datad(\Mux49~15_combout ),
	.cin(gnd),
	.combout(\Mux49~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~16 .lut_mask = 16'hE3E0;
defparam \Mux49~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y41_N25
dffeas \storeregister[5][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][14] .is_wysiwyg = "true";
defparam \storeregister[5][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y41_N19
dffeas \storeregister[4][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][14] .is_wysiwyg = "true";
defparam \storeregister[4][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N24
cycloneive_lcell_comb \Mux49~10 (
// Equation(s):
// \Mux49~10_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][14]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & ((\storeregister[4][14]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][14]~q ),
	.datad(\storeregister[4][14]~q ),
	.cin(gnd),
	.combout(\Mux49~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~10 .lut_mask = 16'hB9A8;
defparam \Mux49~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N18
cycloneive_lcell_comb \Mux49~11 (
// Equation(s):
// \Mux49~11_combout  = (temp_imemload_output_17 & ((\Mux49~10_combout  & (\storeregister[7][14]~q )) # (!\Mux49~10_combout  & ((\storeregister[6][14]~q ))))) # (!temp_imemload_output_17 & (((\Mux49~10_combout ))))

	.dataa(\storeregister[7][14]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[6][14]~q ),
	.datad(\Mux49~10_combout ),
	.cin(gnd),
	.combout(\Mux49~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~11 .lut_mask = 16'hBBC0;
defparam \Mux49~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N8
cycloneive_lcell_comb \Mux54~7 (
// Equation(s):
// \Mux54~7_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[23][9]~q ))) # (!temp_imemload_output_18 & (\storeregister[19][9]~q ))))

	.dataa(\storeregister[19][9]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[23][9]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux54~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~7 .lut_mask = 16'hFC22;
defparam \Mux54~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N26
cycloneive_lcell_comb \Mux54~8 (
// Equation(s):
// \Mux54~8_combout  = (temp_imemload_output_19 & ((\Mux54~7_combout  & (\storeregister[31][9]~q )) # (!\Mux54~7_combout  & ((\storeregister[27][9]~q ))))) # (!temp_imemload_output_19 & (\Mux54~7_combout ))

	.dataa(temp_imemload_output_19),
	.datab(\Mux54~7_combout ),
	.datac(\storeregister[31][9]~q ),
	.datad(\storeregister[27][9]~q ),
	.cin(gnd),
	.combout(\Mux54~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~8 .lut_mask = 16'hE6C4;
defparam \Mux54~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N24
cycloneive_lcell_comb \Mux54~0 (
// Equation(s):
// \Mux54~0_combout  = (temp_imemload_output_18 & ((\storeregister[21][9]~q ) # ((temp_imemload_output_19)))) # (!temp_imemload_output_18 & (((\storeregister[17][9]~q  & !temp_imemload_output_19))))

	.dataa(\storeregister[21][9]~q ),
	.datab(\storeregister[17][9]~q ),
	.datac(temp_imemload_output_18),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~0 .lut_mask = 16'hF0AC;
defparam \Mux54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N12
cycloneive_lcell_comb \storeregister[25][9]~feeder (
// Equation(s):
// \storeregister[25][9]~feeder_combout  = Mux22

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux22),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[25][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[25][9]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[25][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N13
dffeas \storeregister[25][9] (
	.clk(!CLK),
	.d(\storeregister[25][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[25][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[25][9] .is_wysiwyg = "true";
defparam \storeregister[25][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N22
cycloneive_lcell_comb \Mux54~1 (
// Equation(s):
// \Mux54~1_combout  = (temp_imemload_output_19 & ((\Mux54~0_combout  & (\storeregister[29][9]~q )) # (!\Mux54~0_combout  & ((\storeregister[25][9]~q ))))) # (!temp_imemload_output_19 & (\Mux54~0_combout ))

	.dataa(temp_imemload_output_19),
	.datab(\Mux54~0_combout ),
	.datac(\storeregister[29][9]~q ),
	.datad(\storeregister[25][9]~q ),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~1 .lut_mask = 16'hE6C4;
defparam \Mux54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N5
dffeas \storeregister[22][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][9] .is_wysiwyg = "true";
defparam \storeregister[22][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N14
cycloneive_lcell_comb \Mux54~3 (
// Equation(s):
// \Mux54~3_combout  = (\Mux54~2_combout  & (((\storeregister[30][9]~q ) # (!temp_imemload_output_18)))) # (!\Mux54~2_combout  & (\storeregister[22][9]~q  & ((temp_imemload_output_18))))

	.dataa(\Mux54~2_combout ),
	.datab(\storeregister[22][9]~q ),
	.datac(\storeregister[30][9]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux54~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~3 .lut_mask = 16'hE4AA;
defparam \Mux54~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N25
dffeas \storeregister[16][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][9] .is_wysiwyg = "true";
defparam \storeregister[16][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N24
cycloneive_lcell_comb \Mux54~4 (
// Equation(s):
// \Mux54~4_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[24][9]~q ))) # (!temp_imemload_output_19 & (\storeregister[16][9]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[16][9]~q ),
	.datad(\storeregister[24][9]~q ),
	.cin(gnd),
	.combout(\Mux54~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~4 .lut_mask = 16'hDC98;
defparam \Mux54~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N20
cycloneive_lcell_comb \storeregister[20][9]~feeder (
// Equation(s):
// \storeregister[20][9]~feeder_combout  = Mux22

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux22),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[20][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][9]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[20][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N21
dffeas \storeregister[20][9] (
	.clk(!CLK),
	.d(\storeregister[20][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][9] .is_wysiwyg = "true";
defparam \storeregister[20][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N8
cycloneive_lcell_comb \Mux54~5 (
// Equation(s):
// \Mux54~5_combout  = (temp_imemload_output_18 & ((\Mux54~4_combout  & (\storeregister[28][9]~q )) # (!\Mux54~4_combout  & ((\storeregister[20][9]~q ))))) # (!temp_imemload_output_18 & (((\Mux54~4_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[28][9]~q ),
	.datac(\Mux54~4_combout ),
	.datad(\storeregister[20][9]~q ),
	.cin(gnd),
	.combout(\Mux54~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~5 .lut_mask = 16'hDAD0;
defparam \Mux54~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N14
cycloneive_lcell_comb \Mux54~6 (
// Equation(s):
// \Mux54~6_combout  = (temp_imemload_output_17 & ((\Mux54~3_combout ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((\Mux54~5_combout  & !temp_imemload_output_16))))

	.dataa(\Mux54~3_combout ),
	.datab(\Mux54~5_combout ),
	.datac(temp_imemload_output_17),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux54~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~6 .lut_mask = 16'hF0AC;
defparam \Mux54~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N28
cycloneive_lcell_comb \Mux54~17 (
// Equation(s):
// \Mux54~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[13][9]~q )) # (!temp_imemload_output_16 & ((\storeregister[12][9]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[13][9]~q ),
	.datad(\storeregister[12][9]~q ),
	.cin(gnd),
	.combout(\Mux54~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~17 .lut_mask = 16'hD9C8;
defparam \Mux54~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N2
cycloneive_lcell_comb \Mux54~18 (
// Equation(s):
// \Mux54~18_combout  = (\Mux54~17_combout  & (((\storeregister[15][9]~q )) # (!temp_imemload_output_17))) # (!\Mux54~17_combout  & (temp_imemload_output_17 & (\storeregister[14][9]~q )))

	.dataa(\Mux54~17_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[14][9]~q ),
	.datad(\storeregister[15][9]~q ),
	.cin(gnd),
	.combout(\Mux54~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~18 .lut_mask = 16'hEA62;
defparam \Mux54~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y41_N23
dffeas \storeregister[4][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][9] .is_wysiwyg = "true";
defparam \storeregister[4][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N22
cycloneive_lcell_comb \Mux54~12 (
// Equation(s):
// \Mux54~12_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][9]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & (\storeregister[4][9]~q )))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[4][9]~q ),
	.datad(\storeregister[5][9]~q ),
	.cin(gnd),
	.combout(\Mux54~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~12 .lut_mask = 16'hBA98;
defparam \Mux54~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N28
cycloneive_lcell_comb \Mux54~13 (
// Equation(s):
// \Mux54~13_combout  = (temp_imemload_output_17 & ((\Mux54~12_combout  & ((\storeregister[7][9]~q ))) # (!\Mux54~12_combout  & (\storeregister[6][9]~q )))) # (!temp_imemload_output_17 & (((\Mux54~12_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[6][9]~q ),
	.datac(\storeregister[7][9]~q ),
	.datad(\Mux54~12_combout ),
	.cin(gnd),
	.combout(\Mux54~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~13 .lut_mask = 16'hF588;
defparam \Mux54~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N27
dffeas \storeregister[1][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][9] .is_wysiwyg = "true";
defparam \storeregister[1][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N26
cycloneive_lcell_comb \Mux54~14 (
// Equation(s):
// \Mux54~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[3][9]~q ))) # (!temp_imemload_output_17 & (\storeregister[1][9]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[1][9]~q ),
	.datad(\storeregister[3][9]~q ),
	.cin(gnd),
	.combout(\Mux54~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~14 .lut_mask = 16'hC840;
defparam \Mux54~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N14
cycloneive_lcell_comb \Mux54~15 (
// Equation(s):
// \Mux54~15_combout  = (\Mux54~14_combout ) # ((\storeregister[2][9]~q  & (temp_imemload_output_17 & !temp_imemload_output_16)))

	.dataa(\storeregister[2][9]~q ),
	.datab(\Mux54~14_combout ),
	.datac(temp_imemload_output_17),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux54~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~15 .lut_mask = 16'hCCEC;
defparam \Mux54~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N26
cycloneive_lcell_comb \Mux54~16 (
// Equation(s):
// \Mux54~16_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\Mux54~13_combout )) # (!temp_imemload_output_18 & ((\Mux54~15_combout )))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\Mux54~13_combout ),
	.datad(\Mux54~15_combout ),
	.cin(gnd),
	.combout(\Mux54~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~16 .lut_mask = 16'hD9C8;
defparam \Mux54~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N12
cycloneive_lcell_comb \Mux54~10 (
// Equation(s):
// \Mux54~10_combout  = (temp_imemload_output_16 & (temp_imemload_output_17)) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[10][9]~q )) # (!temp_imemload_output_17 & ((\storeregister[8][9]~q )))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[10][9]~q ),
	.datad(\storeregister[8][9]~q ),
	.cin(gnd),
	.combout(\Mux54~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~10 .lut_mask = 16'hD9C8;
defparam \Mux54~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N2
cycloneive_lcell_comb \Mux54~11 (
// Equation(s):
// \Mux54~11_combout  = (\Mux54~10_combout  & (((\storeregister[11][9]~q )) # (!temp_imemload_output_16))) # (!\Mux54~10_combout  & (temp_imemload_output_16 & (\storeregister[9][9]~q )))

	.dataa(\Mux54~10_combout ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[9][9]~q ),
	.datad(\storeregister[11][9]~q ),
	.cin(gnd),
	.combout(\Mux54~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~11 .lut_mask = 16'hEA62;
defparam \Mux54~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N8
cycloneive_lcell_comb \Mux55~7 (
// Equation(s):
// \Mux55~7_combout  = (temp_imemload_output_19 & ((\storeregister[27][8]~q ) # ((temp_imemload_output_18)))) # (!temp_imemload_output_19 & (((\storeregister[19][8]~q  & !temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[27][8]~q ),
	.datac(\storeregister[19][8]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux55~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~7 .lut_mask = 16'hAAD8;
defparam \Mux55~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N26
cycloneive_lcell_comb \Mux55~8 (
// Equation(s):
// \Mux55~8_combout  = (temp_imemload_output_18 & ((\Mux55~7_combout  & (\storeregister[31][8]~q )) # (!\Mux55~7_combout  & ((\storeregister[23][8]~q ))))) # (!temp_imemload_output_18 & (((\Mux55~7_combout ))))

	.dataa(\storeregister[31][8]~q ),
	.datab(\storeregister[23][8]~q ),
	.datac(temp_imemload_output_18),
	.datad(\Mux55~7_combout ),
	.cin(gnd),
	.combout(\Mux55~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~8 .lut_mask = 16'hAFC0;
defparam \Mux55~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N24
cycloneive_lcell_comb \Mux55~0 (
// Equation(s):
// \Mux55~0_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[25][8]~q ))) # (!temp_imemload_output_19 & (\storeregister[17][8]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[17][8]~q ),
	.datad(\storeregister[25][8]~q ),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~0 .lut_mask = 16'hDC98;
defparam \Mux55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N14
cycloneive_lcell_comb \Mux55~1 (
// Equation(s):
// \Mux55~1_combout  = (\Mux55~0_combout  & ((\storeregister[29][8]~q ) # ((!temp_imemload_output_18)))) # (!\Mux55~0_combout  & (((temp_imemload_output_18 & \storeregister[21][8]~q ))))

	.dataa(\storeregister[29][8]~q ),
	.datab(\Mux55~0_combout ),
	.datac(temp_imemload_output_18),
	.datad(\storeregister[21][8]~q ),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~1 .lut_mask = 16'hBC8C;
defparam \Mux55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N17
dffeas \storeregister[22][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][8] .is_wysiwyg = "true";
defparam \storeregister[22][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N16
cycloneive_lcell_comb \Mux55~2 (
// Equation(s):
// \Mux55~2_combout  = (temp_imemload_output_18 & (((\storeregister[22][8]~q ) # (temp_imemload_output_19)))) # (!temp_imemload_output_18 & (\storeregister[18][8]~q  & ((!temp_imemload_output_19))))

	.dataa(\storeregister[18][8]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[22][8]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux55~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~2 .lut_mask = 16'hCCE2;
defparam \Mux55~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N16
cycloneive_lcell_comb \Mux55~3 (
// Equation(s):
// \Mux55~3_combout  = (temp_imemload_output_19 & ((\Mux55~2_combout  & (\storeregister[30][8]~q )) # (!\Mux55~2_combout  & ((\storeregister[26][8]~q ))))) # (!temp_imemload_output_19 & (((\Mux55~2_combout ))))

	.dataa(\storeregister[30][8]~q ),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[26][8]~q ),
	.datad(\Mux55~2_combout ),
	.cin(gnd),
	.combout(\Mux55~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~3 .lut_mask = 16'hBBC0;
defparam \Mux55~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N24
cycloneive_lcell_comb \storeregister[24][8]~feeder (
// Equation(s):
// \storeregister[24][8]~feeder_combout  = Mux23

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux23),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[24][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][8]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[24][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N25
dffeas \storeregister[24][8] (
	.clk(!CLK),
	.d(\storeregister[24][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][8] .is_wysiwyg = "true";
defparam \storeregister[24][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N20
cycloneive_lcell_comb \Mux55~5 (
// Equation(s):
// \Mux55~5_combout  = (\Mux55~4_combout  & (((\storeregister[28][8]~q ) # (!temp_imemload_output_19)))) # (!\Mux55~4_combout  & (\storeregister[24][8]~q  & ((temp_imemload_output_19))))

	.dataa(\Mux55~4_combout ),
	.datab(\storeregister[24][8]~q ),
	.datac(\storeregister[28][8]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux55~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~5 .lut_mask = 16'hE4AA;
defparam \Mux55~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N12
cycloneive_lcell_comb \Mux55~6 (
// Equation(s):
// \Mux55~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\Mux55~3_combout )) # (!temp_imemload_output_17 & ((\Mux55~5_combout )))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux55~3_combout ),
	.datac(\Mux55~5_combout ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux55~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~6 .lut_mask = 16'hEE50;
defparam \Mux55~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N4
cycloneive_lcell_comb \Mux55~17 (
// Equation(s):
// \Mux55~17_combout  = (temp_imemload_output_16 & ((\storeregister[13][8]~q ) # ((temp_imemload_output_17)))) # (!temp_imemload_output_16 & (((\storeregister[12][8]~q  & !temp_imemload_output_17))))

	.dataa(\storeregister[13][8]~q ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[12][8]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux55~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~17 .lut_mask = 16'hCCB8;
defparam \Mux55~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N20
cycloneive_lcell_comb \Mux55~18 (
// Equation(s):
// \Mux55~18_combout  = (temp_imemload_output_17 & ((\Mux55~17_combout  & ((\storeregister[15][8]~q ))) # (!\Mux55~17_combout  & (\storeregister[14][8]~q )))) # (!temp_imemload_output_17 & (((\Mux55~17_combout ))))

	.dataa(\storeregister[14][8]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[15][8]~q ),
	.datad(\Mux55~17_combout ),
	.cin(gnd),
	.combout(\Mux55~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~18 .lut_mask = 16'hF388;
defparam \Mux55~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y41_N1
dffeas \storeregister[5][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][8] .is_wysiwyg = "true";
defparam \storeregister[5][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y41_N11
dffeas \storeregister[4][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][8] .is_wysiwyg = "true";
defparam \storeregister[4][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N0
cycloneive_lcell_comb \Mux55~10 (
// Equation(s):
// \Mux55~10_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][8]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & ((\storeregister[4][8]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[5][8]~q ),
	.datad(\storeregister[4][8]~q ),
	.cin(gnd),
	.combout(\Mux55~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~10 .lut_mask = 16'hB9A8;
defparam \Mux55~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N28
cycloneive_lcell_comb \Mux55~11 (
// Equation(s):
// \Mux55~11_combout  = (\Mux55~10_combout  & ((\storeregister[7][8]~q ) # ((!temp_imemload_output_17)))) # (!\Mux55~10_combout  & (((\storeregister[6][8]~q  & temp_imemload_output_17))))

	.dataa(\storeregister[7][8]~q ),
	.datab(\Mux55~10_combout ),
	.datac(\storeregister[6][8]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux55~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~11 .lut_mask = 16'hB8CC;
defparam \Mux55~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N4
cycloneive_lcell_comb \Mux55~12 (
// Equation(s):
// \Mux55~12_combout  = (temp_imemload_output_16 & (temp_imemload_output_17)) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[10][8]~q ))) # (!temp_imemload_output_17 & (\storeregister[8][8]~q ))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[8][8]~q ),
	.datad(\storeregister[10][8]~q ),
	.cin(gnd),
	.combout(\Mux55~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~12 .lut_mask = 16'hDC98;
defparam \Mux55~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N6
cycloneive_lcell_comb \Mux55~13 (
// Equation(s):
// \Mux55~13_combout  = (temp_imemload_output_16 & ((\Mux55~12_combout  & (\storeregister[11][8]~q )) # (!\Mux55~12_combout  & ((\storeregister[9][8]~q ))))) # (!temp_imemload_output_16 & (\Mux55~12_combout ))

	.dataa(temp_imemload_output_16),
	.datab(\Mux55~12_combout ),
	.datac(\storeregister[11][8]~q ),
	.datad(\storeregister[9][8]~q ),
	.cin(gnd),
	.combout(\Mux55~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~13 .lut_mask = 16'hE6C4;
defparam \Mux55~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N13
dffeas \storeregister[3][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[3][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[3][8] .is_wysiwyg = "true";
defparam \storeregister[3][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N3
dffeas \storeregister[1][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[1][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[1][8] .is_wysiwyg = "true";
defparam \storeregister[1][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N12
cycloneive_lcell_comb \Mux55~14 (
// Equation(s):
// \Mux55~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][8]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][8]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[3][8]~q ),
	.datad(\storeregister[1][8]~q ),
	.cin(gnd),
	.combout(\Mux55~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~14 .lut_mask = 16'hC480;
defparam \Mux55~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N10
cycloneive_lcell_comb \Mux55~15 (
// Equation(s):
// \Mux55~15_combout  = (\Mux55~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][8]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux55~14_combout ),
	.datac(\storeregister[2][8]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux55~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~15 .lut_mask = 16'hCCEC;
defparam \Mux55~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N10
cycloneive_lcell_comb \Mux55~16 (
// Equation(s):
// \Mux55~16_combout  = (temp_imemload_output_19 & ((temp_imemload_output_18) # ((\Mux55~13_combout )))) # (!temp_imemload_output_19 & (!temp_imemload_output_18 & ((\Mux55~15_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\Mux55~13_combout ),
	.datad(\Mux55~15_combout ),
	.cin(gnd),
	.combout(\Mux55~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~16 .lut_mask = 16'hB9A8;
defparam \Mux55~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N26
cycloneive_lcell_comb \Mux56~0 (
// Equation(s):
// \Mux56~0_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[21][7]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[17][7]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[21][7]~q ),
	.datad(\storeregister[17][7]~q ),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~0 .lut_mask = 16'hB9A8;
defparam \Mux56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N12
cycloneive_lcell_comb \Mux56~1 (
// Equation(s):
// \Mux56~1_combout  = (\Mux56~0_combout  & ((\storeregister[29][7]~q ) # ((!temp_imemload_output_19)))) # (!\Mux56~0_combout  & (((temp_imemload_output_19 & \storeregister[25][7]~q ))))

	.dataa(\Mux56~0_combout ),
	.datab(\storeregister[29][7]~q ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[25][7]~q ),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~1 .lut_mask = 16'hDA8A;
defparam \Mux56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N2
cycloneive_lcell_comb \Mux56~7 (
// Equation(s):
// \Mux56~7_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[23][7]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[19][7]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[19][7]~q ),
	.datad(\storeregister[23][7]~q ),
	.cin(gnd),
	.combout(\Mux56~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~7 .lut_mask = 16'hBA98;
defparam \Mux56~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N4
cycloneive_lcell_comb \Mux56~8 (
// Equation(s):
// \Mux56~8_combout  = (temp_imemload_output_19 & ((\Mux56~7_combout  & (\storeregister[31][7]~q )) # (!\Mux56~7_combout  & ((\storeregister[27][7]~q ))))) # (!temp_imemload_output_19 & (((\Mux56~7_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[31][7]~q ),
	.datac(\storeregister[27][7]~q ),
	.datad(\Mux56~7_combout ),
	.cin(gnd),
	.combout(\Mux56~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~8 .lut_mask = 16'hDDA0;
defparam \Mux56~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N22
cycloneive_lcell_comb \Mux56~4 (
// Equation(s):
// \Mux56~4_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[24][7]~q ))) # (!temp_imemload_output_19 & (\storeregister[16][7]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[16][7]~q ),
	.datad(\storeregister[24][7]~q ),
	.cin(gnd),
	.combout(\Mux56~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~4 .lut_mask = 16'hDC98;
defparam \Mux56~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N30
cycloneive_lcell_comb \Mux56~5 (
// Equation(s):
// \Mux56~5_combout  = (temp_imemload_output_18 & ((\Mux56~4_combout  & (\storeregister[28][7]~q )) # (!\Mux56~4_combout  & ((\storeregister[20][7]~q ))))) # (!temp_imemload_output_18 & (\Mux56~4_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux56~4_combout ),
	.datac(\storeregister[28][7]~q ),
	.datad(\storeregister[20][7]~q ),
	.cin(gnd),
	.combout(\Mux56~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~5 .lut_mask = 16'hE6C4;
defparam \Mux56~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N22
cycloneive_lcell_comb \Mux56~3 (
// Equation(s):
// \Mux56~3_combout  = (\Mux56~2_combout  & ((\storeregister[30][7]~q ) # ((!temp_imemload_output_18)))) # (!\Mux56~2_combout  & (((\storeregister[22][7]~q  & temp_imemload_output_18))))

	.dataa(\Mux56~2_combout ),
	.datab(\storeregister[30][7]~q ),
	.datac(\storeregister[22][7]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux56~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~3 .lut_mask = 16'hD8AA;
defparam \Mux56~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N26
cycloneive_lcell_comb \Mux56~6 (
// Equation(s):
// \Mux56~6_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16) # (\Mux56~3_combout )))) # (!temp_imemload_output_17 & (\Mux56~5_combout  & (!temp_imemload_output_16)))

	.dataa(\Mux56~5_combout ),
	.datab(temp_imemload_output_17),
	.datac(temp_imemload_output_16),
	.datad(\Mux56~3_combout ),
	.cin(gnd),
	.combout(\Mux56~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~6 .lut_mask = 16'hCEC2;
defparam \Mux56~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N0
cycloneive_lcell_comb \Mux56~17 (
// Equation(s):
// \Mux56~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][7]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][7]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[12][7]~q ),
	.datad(\storeregister[13][7]~q ),
	.cin(gnd),
	.combout(\Mux56~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~17 .lut_mask = 16'hDC98;
defparam \Mux56~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N20
cycloneive_lcell_comb \Mux56~18 (
// Equation(s):
// \Mux56~18_combout  = (temp_imemload_output_17 & ((\Mux56~17_combout  & ((\storeregister[15][7]~q ))) # (!\Mux56~17_combout  & (\storeregister[14][7]~q )))) # (!temp_imemload_output_17 & (((\Mux56~17_combout ))))

	.dataa(\storeregister[14][7]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[15][7]~q ),
	.datad(\Mux56~17_combout ),
	.cin(gnd),
	.combout(\Mux56~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~18 .lut_mask = 16'hF388;
defparam \Mux56~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N4
cycloneive_lcell_comb \Mux56~14 (
// Equation(s):
// \Mux56~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][7]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][7]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[3][7]~q ),
	.datad(\storeregister[1][7]~q ),
	.cin(gnd),
	.combout(\Mux56~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~14 .lut_mask = 16'hC480;
defparam \Mux56~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N26
cycloneive_lcell_comb \Mux56~15 (
// Equation(s):
// \Mux56~15_combout  = (\Mux56~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][7]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux56~14_combout ),
	.datac(\storeregister[2][7]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux56~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~15 .lut_mask = 16'hCCEC;
defparam \Mux56~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N4
cycloneive_lcell_comb \Mux56~13 (
// Equation(s):
// \Mux56~13_combout  = (\Mux56~12_combout  & (((\storeregister[7][7]~q )) # (!temp_imemload_output_17))) # (!\Mux56~12_combout  & (temp_imemload_output_17 & (\storeregister[6][7]~q )))

	.dataa(\Mux56~12_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[6][7]~q ),
	.datad(\storeregister[7][7]~q ),
	.cin(gnd),
	.combout(\Mux56~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~13 .lut_mask = 16'hEA62;
defparam \Mux56~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N8
cycloneive_lcell_comb \Mux56~16 (
// Equation(s):
// \Mux56~16_combout  = (temp_imemload_output_19 & (temp_imemload_output_18)) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\Mux56~13_combout ))) # (!temp_imemload_output_18 & (\Mux56~15_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(temp_imemload_output_18),
	.datac(\Mux56~15_combout ),
	.datad(\Mux56~13_combout ),
	.cin(gnd),
	.combout(\Mux56~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~16 .lut_mask = 16'hDC98;
defparam \Mux56~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N10
cycloneive_lcell_comb \storeregister[11][7]~feeder (
// Equation(s):
// \storeregister[11][7]~feeder_combout  = Mux24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux24),
	.cin(gnd),
	.combout(\storeregister[11][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[11][7]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[11][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N11
dffeas \storeregister[11][7] (
	.clk(!CLK),
	.d(\storeregister[11][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[11][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[11][7] .is_wysiwyg = "true";
defparam \storeregister[11][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N20
cycloneive_lcell_comb \Mux56~10 (
// Equation(s):
// \Mux56~10_combout  = (temp_imemload_output_16 & (temp_imemload_output_17)) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[10][7]~q )) # (!temp_imemload_output_17 & ((\storeregister[8][7]~q )))))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[10][7]~q ),
	.datad(\storeregister[8][7]~q ),
	.cin(gnd),
	.combout(\Mux56~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~10 .lut_mask = 16'hD9C8;
defparam \Mux56~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N18
cycloneive_lcell_comb \Mux56~11 (
// Equation(s):
// \Mux56~11_combout  = (temp_imemload_output_16 & ((\Mux56~10_combout  & (\storeregister[11][7]~q )) # (!\Mux56~10_combout  & ((\storeregister[9][7]~q ))))) # (!temp_imemload_output_16 & (((\Mux56~10_combout ))))

	.dataa(\storeregister[11][7]~q ),
	.datab(temp_imemload_output_16),
	.datac(\Mux56~10_combout ),
	.datad(\storeregister[9][7]~q ),
	.cin(gnd),
	.combout(\Mux56~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~11 .lut_mask = 16'hBCB0;
defparam \Mux56~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N26
cycloneive_lcell_comb \Mux57~7 (
// Equation(s):
// \Mux57~7_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\storeregister[27][6]~q )) # (!temp_imemload_output_19 & ((\storeregister[19][6]~q )))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[27][6]~q ),
	.datad(\storeregister[19][6]~q ),
	.cin(gnd),
	.combout(\Mux57~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~7 .lut_mask = 16'hD9C8;
defparam \Mux57~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N20
cycloneive_lcell_comb \Mux57~8 (
// Equation(s):
// \Mux57~8_combout  = (temp_imemload_output_18 & ((\Mux57~7_combout  & ((\storeregister[31][6]~q ))) # (!\Mux57~7_combout  & (\storeregister[23][6]~q )))) # (!temp_imemload_output_18 & (((\Mux57~7_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[23][6]~q ),
	.datac(\Mux57~7_combout ),
	.datad(\storeregister[31][6]~q ),
	.cin(gnd),
	.combout(\Mux57~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~8 .lut_mask = 16'hF858;
defparam \Mux57~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N28
cycloneive_lcell_comb \Mux57~2 (
// Equation(s):
// \Mux57~2_combout  = (temp_imemload_output_18 & (((\storeregister[22][6]~q ) # (temp_imemload_output_19)))) # (!temp_imemload_output_18 & (\storeregister[18][6]~q  & ((!temp_imemload_output_19))))

	.dataa(\storeregister[18][6]~q ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[22][6]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux57~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~2 .lut_mask = 16'hCCE2;
defparam \Mux57~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N0
cycloneive_lcell_comb \Mux57~3 (
// Equation(s):
// \Mux57~3_combout  = (temp_imemload_output_19 & ((\Mux57~2_combout  & ((\storeregister[30][6]~q ))) # (!\Mux57~2_combout  & (\storeregister[26][6]~q )))) # (!temp_imemload_output_19 & (\Mux57~2_combout ))

	.dataa(temp_imemload_output_19),
	.datab(\Mux57~2_combout ),
	.datac(\storeregister[26][6]~q ),
	.datad(\storeregister[30][6]~q ),
	.cin(gnd),
	.combout(\Mux57~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~3 .lut_mask = 16'hEC64;
defparam \Mux57~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N8
cycloneive_lcell_comb \Mux57~5 (
// Equation(s):
// \Mux57~5_combout  = (\Mux57~4_combout  & ((\storeregister[28][6]~q ) # ((!temp_imemload_output_19)))) # (!\Mux57~4_combout  & (((temp_imemload_output_19 & \storeregister[24][6]~q ))))

	.dataa(\Mux57~4_combout ),
	.datab(\storeregister[28][6]~q ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[24][6]~q ),
	.cin(gnd),
	.combout(\Mux57~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~5 .lut_mask = 16'hDA8A;
defparam \Mux57~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N4
cycloneive_lcell_comb \Mux57~6 (
// Equation(s):
// \Mux57~6_combout  = (temp_imemload_output_17 & ((temp_imemload_output_16) # ((\Mux57~3_combout )))) # (!temp_imemload_output_17 & (!temp_imemload_output_16 & ((\Mux57~5_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\Mux57~3_combout ),
	.datad(\Mux57~5_combout ),
	.cin(gnd),
	.combout(\Mux57~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~6 .lut_mask = 16'hB9A8;
defparam \Mux57~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N13
dffeas \storeregister[17][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][6] .is_wysiwyg = "true";
defparam \storeregister[17][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N12
cycloneive_lcell_comb \Mux57~0 (
// Equation(s):
// \Mux57~0_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[25][6]~q ))) # (!temp_imemload_output_19 & (\storeregister[17][6]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[17][6]~q ),
	.datad(\storeregister[25][6]~q ),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~0 .lut_mask = 16'hDC98;
defparam \Mux57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N10
cycloneive_lcell_comb \Mux57~1 (
// Equation(s):
// \Mux57~1_combout  = (temp_imemload_output_18 & ((\Mux57~0_combout  & ((\storeregister[29][6]~q ))) # (!\Mux57~0_combout  & (\storeregister[21][6]~q )))) # (!temp_imemload_output_18 & (((\Mux57~0_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[21][6]~q ),
	.datac(\Mux57~0_combout ),
	.datad(\storeregister[29][6]~q ),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~1 .lut_mask = 16'hF858;
defparam \Mux57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N28
cycloneive_lcell_comb \Mux57~12 (
// Equation(s):
// \Mux57~12_combout  = (temp_imemload_output_17 & ((\storeregister[10][6]~q ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((\storeregister[8][6]~q  & !temp_imemload_output_16))))

	.dataa(\storeregister[10][6]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[8][6]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux57~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~12 .lut_mask = 16'hCCB8;
defparam \Mux57~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N26
cycloneive_lcell_comb \Mux57~13 (
// Equation(s):
// \Mux57~13_combout  = (temp_imemload_output_16 & ((\Mux57~12_combout  & (\storeregister[11][6]~q )) # (!\Mux57~12_combout  & ((\storeregister[9][6]~q ))))) # (!temp_imemload_output_16 & (\Mux57~12_combout ))

	.dataa(temp_imemload_output_16),
	.datab(\Mux57~12_combout ),
	.datac(\storeregister[11][6]~q ),
	.datad(\storeregister[9][6]~q ),
	.cin(gnd),
	.combout(\Mux57~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~13 .lut_mask = 16'hE6C4;
defparam \Mux57~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N24
cycloneive_lcell_comb \Mux57~14 (
// Equation(s):
// \Mux57~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & (\storeregister[3][6]~q )) # (!temp_imemload_output_17 & ((\storeregister[1][6]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[3][6]~q ),
	.datad(\storeregister[1][6]~q ),
	.cin(gnd),
	.combout(\Mux57~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~14 .lut_mask = 16'hC480;
defparam \Mux57~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N30
cycloneive_lcell_comb \Mux57~15 (
// Equation(s):
// \Mux57~15_combout  = (\Mux57~14_combout ) # ((temp_imemload_output_17 & (!temp_imemload_output_16 & \storeregister[2][6]~q )))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[2][6]~q ),
	.datad(\Mux57~14_combout ),
	.cin(gnd),
	.combout(\Mux57~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~15 .lut_mask = 16'hFF20;
defparam \Mux57~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N6
cycloneive_lcell_comb \Mux57~16 (
// Equation(s):
// \Mux57~16_combout  = (temp_imemload_output_18 & (((temp_imemload_output_19)))) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\Mux57~13_combout )) # (!temp_imemload_output_19 & ((\Mux57~15_combout )))))

	.dataa(\Mux57~13_combout ),
	.datab(temp_imemload_output_18),
	.datac(temp_imemload_output_19),
	.datad(\Mux57~15_combout ),
	.cin(gnd),
	.combout(\Mux57~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~16 .lut_mask = 16'hE3E0;
defparam \Mux57~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y41_N15
dffeas \storeregister[4][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][6] .is_wysiwyg = "true";
defparam \storeregister[4][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y41_N5
dffeas \storeregister[5][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[5][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[5][6] .is_wysiwyg = "true";
defparam \storeregister[5][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N4
cycloneive_lcell_comb \Mux57~10 (
// Equation(s):
// \Mux57~10_combout  = (temp_imemload_output_16 & (((\storeregister[5][6]~q ) # (temp_imemload_output_17)))) # (!temp_imemload_output_16 & (\storeregister[4][6]~q  & ((!temp_imemload_output_17))))

	.dataa(temp_imemload_output_16),
	.datab(\storeregister[4][6]~q ),
	.datac(\storeregister[5][6]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux57~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~10 .lut_mask = 16'hAAE4;
defparam \Mux57~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N24
cycloneive_lcell_comb \Mux57~11 (
// Equation(s):
// \Mux57~11_combout  = (\Mux57~10_combout  & ((\storeregister[7][6]~q ) # ((!temp_imemload_output_17)))) # (!\Mux57~10_combout  & (((\storeregister[6][6]~q  & temp_imemload_output_17))))

	.dataa(\Mux57~10_combout ),
	.datab(\storeregister[7][6]~q ),
	.datac(\storeregister[6][6]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux57~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~11 .lut_mask = 16'hD8AA;
defparam \Mux57~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N16
cycloneive_lcell_comb \Mux57~17 (
// Equation(s):
// \Mux57~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][6]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][6]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[12][6]~q ),
	.datad(\storeregister[13][6]~q ),
	.cin(gnd),
	.combout(\Mux57~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~17 .lut_mask = 16'hDC98;
defparam \Mux57~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N10
cycloneive_lcell_comb \Mux57~18 (
// Equation(s):
// \Mux57~18_combout  = (\Mux57~17_combout  & ((\storeregister[15][6]~q ) # ((!temp_imemload_output_17)))) # (!\Mux57~17_combout  & (((\storeregister[14][6]~q  & temp_imemload_output_17))))

	.dataa(\storeregister[15][6]~q ),
	.datab(\Mux57~17_combout ),
	.datac(\storeregister[14][6]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux57~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~18 .lut_mask = 16'hB8CC;
defparam \Mux57~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N10
cycloneive_lcell_comb \Mux58~0 (
// Equation(s):
// \Mux58~0_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\storeregister[21][5]~q ))) # (!temp_imemload_output_18 & (\storeregister[17][5]~q ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[17][5]~q ),
	.datac(temp_imemload_output_18),
	.datad(\storeregister[21][5]~q ),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~0 .lut_mask = 16'hF4A4;
defparam \Mux58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N8
cycloneive_lcell_comb \Mux58~1 (
// Equation(s):
// \Mux58~1_combout  = (temp_imemload_output_19 & ((\Mux58~0_combout  & (\storeregister[29][5]~q )) # (!\Mux58~0_combout  & ((\storeregister[25][5]~q ))))) # (!temp_imemload_output_19 & (((\Mux58~0_combout ))))

	.dataa(\storeregister[29][5]~q ),
	.datab(\storeregister[25][5]~q ),
	.datac(temp_imemload_output_19),
	.datad(\Mux58~0_combout ),
	.cin(gnd),
	.combout(\Mux58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~1 .lut_mask = 16'hAFC0;
defparam \Mux58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N30
cycloneive_lcell_comb \Mux58~7 (
// Equation(s):
// \Mux58~7_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[23][5]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[19][5]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[19][5]~q ),
	.datad(\storeregister[23][5]~q ),
	.cin(gnd),
	.combout(\Mux58~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~7 .lut_mask = 16'hBA98;
defparam \Mux58~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N14
cycloneive_lcell_comb \Mux58~8 (
// Equation(s):
// \Mux58~8_combout  = (\Mux58~7_combout  & (((\storeregister[31][5]~q ) # (!temp_imemload_output_19)))) # (!\Mux58~7_combout  & (\storeregister[27][5]~q  & ((temp_imemload_output_19))))

	.dataa(\Mux58~7_combout ),
	.datab(\storeregister[27][5]~q ),
	.datac(\storeregister[31][5]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux58~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~8 .lut_mask = 16'hE4AA;
defparam \Mux58~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N5
dffeas \storeregister[16][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][5] .is_wysiwyg = "true";
defparam \storeregister[16][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N2
cycloneive_lcell_comb \storeregister[24][5]~feeder (
// Equation(s):
// \storeregister[24][5]~feeder_combout  = Mux26

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux26),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[24][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[24][5]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[24][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N3
dffeas \storeregister[24][5] (
	.clk(!CLK),
	.d(\storeregister[24][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][5] .is_wysiwyg = "true";
defparam \storeregister[24][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N4
cycloneive_lcell_comb \Mux58~4 (
// Equation(s):
// \Mux58~4_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & ((\storeregister[24][5]~q ))) # (!temp_imemload_output_19 & (\storeregister[16][5]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[16][5]~q ),
	.datad(\storeregister[24][5]~q ),
	.cin(gnd),
	.combout(\Mux58~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~4 .lut_mask = 16'hDC98;
defparam \Mux58~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N26
cycloneive_lcell_comb \Mux58~5 (
// Equation(s):
// \Mux58~5_combout  = (temp_imemload_output_18 & ((\Mux58~4_combout  & (\storeregister[28][5]~q )) # (!\Mux58~4_combout  & ((\storeregister[20][5]~q ))))) # (!temp_imemload_output_18 & (((\Mux58~4_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[28][5]~q ),
	.datac(\Mux58~4_combout ),
	.datad(\storeregister[20][5]~q ),
	.cin(gnd),
	.combout(\Mux58~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~5 .lut_mask = 16'hDAD0;
defparam \Mux58~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N8
cycloneive_lcell_comb \storeregister[22][5]~feeder (
// Equation(s):
// \storeregister[22][5]~feeder_combout  = Mux26

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux26),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[22][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[22][5]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[22][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N9
dffeas \storeregister[22][5] (
	.clk(!CLK),
	.d(\storeregister[22][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[22][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[22][5] .is_wysiwyg = "true";
defparam \storeregister[22][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N7
dffeas \storeregister[30][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[30][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[30][5] .is_wysiwyg = "true";
defparam \storeregister[30][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N6
cycloneive_lcell_comb \Mux58~3 (
// Equation(s):
// \Mux58~3_combout  = (\Mux58~2_combout  & (((\storeregister[30][5]~q ) # (!temp_imemload_output_18)))) # (!\Mux58~2_combout  & (\storeregister[22][5]~q  & ((temp_imemload_output_18))))

	.dataa(\Mux58~2_combout ),
	.datab(\storeregister[22][5]~q ),
	.datac(\storeregister[30][5]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux58~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~3 .lut_mask = 16'hE4AA;
defparam \Mux58~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N16
cycloneive_lcell_comb \Mux58~6 (
// Equation(s):
// \Mux58~6_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16) # (\Mux58~3_combout )))) # (!temp_imemload_output_17 & (\Mux58~5_combout  & (!temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux58~5_combout ),
	.datac(temp_imemload_output_16),
	.datad(\Mux58~3_combout ),
	.cin(gnd),
	.combout(\Mux58~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~6 .lut_mask = 16'hAEA4;
defparam \Mux58~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N12
cycloneive_lcell_comb \Mux58~17 (
// Equation(s):
// \Mux58~17_combout  = (temp_imemload_output_17 & (temp_imemload_output_16)) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][5]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][5]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[12][5]~q ),
	.datad(\storeregister[13][5]~q ),
	.cin(gnd),
	.combout(\Mux58~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~17 .lut_mask = 16'hDC98;
defparam \Mux58~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N26
cycloneive_lcell_comb \Mux58~18 (
// Equation(s):
// \Mux58~18_combout  = (temp_imemload_output_17 & ((\Mux58~17_combout  & (\storeregister[15][5]~q )) # (!\Mux58~17_combout  & ((\storeregister[14][5]~q ))))) # (!temp_imemload_output_17 & (((\Mux58~17_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[15][5]~q ),
	.datac(\storeregister[14][5]~q ),
	.datad(\Mux58~17_combout ),
	.cin(gnd),
	.combout(\Mux58~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~18 .lut_mask = 16'hDDA0;
defparam \Mux58~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N25
dffeas \storeregister[10][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][5] .is_wysiwyg = "true";
defparam \storeregister[10][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N24
cycloneive_lcell_comb \Mux58~10 (
// Equation(s):
// \Mux58~10_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[10][5]~q ))) # (!temp_imemload_output_17 & (\storeregister[8][5]~q ))))

	.dataa(\storeregister[8][5]~q ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[10][5]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux58~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~10 .lut_mask = 16'hFC22;
defparam \Mux58~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N28
cycloneive_lcell_comb \Mux58~11 (
// Equation(s):
// \Mux58~11_combout  = (\Mux58~10_combout  & ((\storeregister[11][5]~q ) # ((!temp_imemload_output_16)))) # (!\Mux58~10_combout  & (((\storeregister[9][5]~q  & temp_imemload_output_16))))

	.dataa(\storeregister[11][5]~q ),
	.datab(\Mux58~10_combout ),
	.datac(\storeregister[9][5]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux58~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~11 .lut_mask = 16'hB8CC;
defparam \Mux58~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N26
cycloneive_lcell_comb \Mux58~12 (
// Equation(s):
// \Mux58~12_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][5]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & (\storeregister[4][5]~q )))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[4][5]~q ),
	.datad(\storeregister[5][5]~q ),
	.cin(gnd),
	.combout(\Mux58~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~12 .lut_mask = 16'hBA98;
defparam \Mux58~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N16
cycloneive_lcell_comb \Mux58~13 (
// Equation(s):
// \Mux58~13_combout  = (temp_imemload_output_17 & ((\Mux58~12_combout  & ((\storeregister[7][5]~q ))) # (!\Mux58~12_combout  & (\storeregister[6][5]~q )))) # (!temp_imemload_output_17 & (((\Mux58~12_combout ))))

	.dataa(\storeregister[6][5]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[7][5]~q ),
	.datad(\Mux58~12_combout ),
	.cin(gnd),
	.combout(\Mux58~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~13 .lut_mask = 16'hF388;
defparam \Mux58~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N28
cycloneive_lcell_comb \Mux58~14 (
// Equation(s):
// \Mux58~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[3][5]~q ))) # (!temp_imemload_output_17 & (\storeregister[1][5]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[1][5]~q ),
	.datac(\storeregister[3][5]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux58~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~14 .lut_mask = 16'hE400;
defparam \Mux58~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N14
cycloneive_lcell_comb \Mux58~15 (
// Equation(s):
// \Mux58~15_combout  = (\Mux58~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][5]~q  & !temp_imemload_output_16)))

	.dataa(temp_imemload_output_17),
	.datab(\Mux58~14_combout ),
	.datac(\storeregister[2][5]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux58~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~15 .lut_mask = 16'hCCEC;
defparam \Mux58~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N28
cycloneive_lcell_comb \Mux58~16 (
// Equation(s):
// \Mux58~16_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & (\Mux58~13_combout )) # (!temp_imemload_output_18 & ((\Mux58~15_combout )))))

	.dataa(temp_imemload_output_19),
	.datab(\Mux58~13_combout ),
	.datac(\Mux58~15_combout ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux58~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~16 .lut_mask = 16'hEE50;
defparam \Mux58~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N16
cycloneive_lcell_comb \Mux50~7 (
// Equation(s):
// \Mux50~7_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[23][13]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\storeregister[19][13]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[23][13]~q ),
	.datad(\storeregister[19][13]~q ),
	.cin(gnd),
	.combout(\Mux50~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~7 .lut_mask = 16'hB9A8;
defparam \Mux50~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N20
cycloneive_lcell_comb \Mux50~8 (
// Equation(s):
// \Mux50~8_combout  = (temp_imemload_output_19 & ((\Mux50~7_combout  & (\storeregister[31][13]~q )) # (!\Mux50~7_combout  & ((\storeregister[27][13]~q ))))) # (!temp_imemload_output_19 & (((\Mux50~7_combout ))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[31][13]~q ),
	.datac(\storeregister[27][13]~q ),
	.datad(\Mux50~7_combout ),
	.cin(gnd),
	.combout(\Mux50~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~8 .lut_mask = 16'hDDA0;
defparam \Mux50~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N16
cycloneive_lcell_comb \Mux50~3 (
// Equation(s):
// \Mux50~3_combout  = (\Mux50~2_combout  & (((\storeregister[30][13]~q )) # (!temp_imemload_output_18))) # (!\Mux50~2_combout  & (temp_imemload_output_18 & (\storeregister[22][13]~q )))

	.dataa(\Mux50~2_combout ),
	.datab(temp_imemload_output_18),
	.datac(\storeregister[22][13]~q ),
	.datad(\storeregister[30][13]~q ),
	.cin(gnd),
	.combout(\Mux50~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~3 .lut_mask = 16'hEA62;
defparam \Mux50~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N28
cycloneive_lcell_comb \storeregister[16][13]~feeder (
// Equation(s):
// \storeregister[16][13]~feeder_combout  = Mux18

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux18),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[16][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[16][13]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[16][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N29
dffeas \storeregister[16][13] (
	.clk(!CLK),
	.d(\storeregister[16][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[16][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[16][13] .is_wysiwyg = "true";
defparam \storeregister[16][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N18
cycloneive_lcell_comb \Mux50~4 (
// Equation(s):
// \Mux50~4_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\storeregister[24][13]~q )) # (!temp_imemload_output_19 & ((\storeregister[16][13]~q )))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[24][13]~q ),
	.datad(\storeregister[16][13]~q ),
	.cin(gnd),
	.combout(\Mux50~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~4 .lut_mask = 16'hD9C8;
defparam \Mux50~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N18
cycloneive_lcell_comb \Mux50~5 (
// Equation(s):
// \Mux50~5_combout  = (temp_imemload_output_18 & ((\Mux50~4_combout  & ((\storeregister[28][13]~q ))) # (!\Mux50~4_combout  & (\storeregister[20][13]~q )))) # (!temp_imemload_output_18 & (((\Mux50~4_combout ))))

	.dataa(\storeregister[20][13]~q ),
	.datab(\storeregister[28][13]~q ),
	.datac(temp_imemload_output_18),
	.datad(\Mux50~4_combout ),
	.cin(gnd),
	.combout(\Mux50~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~5 .lut_mask = 16'hCFA0;
defparam \Mux50~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N8
cycloneive_lcell_comb \Mux50~6 (
// Equation(s):
// \Mux50~6_combout  = (temp_imemload_output_17 & ((\Mux50~3_combout ) # ((temp_imemload_output_16)))) # (!temp_imemload_output_17 & (((\Mux50~5_combout  & !temp_imemload_output_16))))

	.dataa(\Mux50~3_combout ),
	.datab(\Mux50~5_combout ),
	.datac(temp_imemload_output_17),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux50~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~6 .lut_mask = 16'hF0AC;
defparam \Mux50~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N15
dffeas \storeregister[17][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[17][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[17][13] .is_wysiwyg = "true";
defparam \storeregister[17][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N14
cycloneive_lcell_comb \Mux50~0 (
// Equation(s):
// \Mux50~0_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\storeregister[21][13]~q )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & (\storeregister[17][13]~q )))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[17][13]~q ),
	.datad(\storeregister[21][13]~q ),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~0 .lut_mask = 16'hBA98;
defparam \Mux50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N26
cycloneive_lcell_comb \Mux50~1 (
// Equation(s):
// \Mux50~1_combout  = (\Mux50~0_combout  & (((\storeregister[29][13]~q ) # (!temp_imemload_output_19)))) # (!\Mux50~0_combout  & (\storeregister[25][13]~q  & (temp_imemload_output_19)))

	.dataa(\Mux50~0_combout ),
	.datab(\storeregister[25][13]~q ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[29][13]~q ),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~1 .lut_mask = 16'hEA4A;
defparam \Mux50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N5
dffeas \storeregister[10][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][13] .is_wysiwyg = "true";
defparam \storeregister[10][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N4
cycloneive_lcell_comb \Mux50~10 (
// Equation(s):
// \Mux50~10_combout  = (temp_imemload_output_17 & (((\storeregister[10][13]~q ) # (temp_imemload_output_16)))) # (!temp_imemload_output_17 & (\storeregister[8][13]~q  & ((!temp_imemload_output_16))))

	.dataa(\storeregister[8][13]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[10][13]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux50~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~10 .lut_mask = 16'hCCE2;
defparam \Mux50~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N12
cycloneive_lcell_comb \Mux50~11 (
// Equation(s):
// \Mux50~11_combout  = (\Mux50~10_combout  & ((\storeregister[11][13]~q ) # ((!temp_imemload_output_16)))) # (!\Mux50~10_combout  & (((\storeregister[9][13]~q  & temp_imemload_output_16))))

	.dataa(\storeregister[11][13]~q ),
	.datab(\Mux50~10_combout ),
	.datac(\storeregister[9][13]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux50~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~11 .lut_mask = 16'hB8CC;
defparam \Mux50~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N22
cycloneive_lcell_comb \Mux50~14 (
// Equation(s):
// \Mux50~14_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17 & ((\storeregister[3][13]~q ))) # (!temp_imemload_output_17 & (\storeregister[1][13]~q ))))

	.dataa(temp_imemload_output_17),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[1][13]~q ),
	.datad(\storeregister[3][13]~q ),
	.cin(gnd),
	.combout(\Mux50~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~14 .lut_mask = 16'hC840;
defparam \Mux50~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N22
cycloneive_lcell_comb \Mux50~15 (
// Equation(s):
// \Mux50~15_combout  = (\Mux50~14_combout ) # ((!temp_imemload_output_16 & (temp_imemload_output_17 & \storeregister[2][13]~q )))

	.dataa(temp_imemload_output_16),
	.datab(\Mux50~14_combout ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[2][13]~q ),
	.cin(gnd),
	.combout(\Mux50~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~15 .lut_mask = 16'hDCCC;
defparam \Mux50~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y41_N31
dffeas \storeregister[4][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[4][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[4][13] .is_wysiwyg = "true";
defparam \storeregister[4][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y41_N30
cycloneive_lcell_comb \Mux50~12 (
// Equation(s):
// \Mux50~12_combout  = (temp_imemload_output_16 & ((temp_imemload_output_17) # ((\storeregister[5][13]~q )))) # (!temp_imemload_output_16 & (!temp_imemload_output_17 & (\storeregister[4][13]~q )))

	.dataa(temp_imemload_output_16),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[4][13]~q ),
	.datad(\storeregister[5][13]~q ),
	.cin(gnd),
	.combout(\Mux50~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~12 .lut_mask = 16'hBA98;
defparam \Mux50~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y39_N6
cycloneive_lcell_comb \Mux50~13 (
// Equation(s):
// \Mux50~13_combout  = (temp_imemload_output_17 & ((\Mux50~12_combout  & ((\storeregister[7][13]~q ))) # (!\Mux50~12_combout  & (\storeregister[6][13]~q )))) # (!temp_imemload_output_17 & (((\Mux50~12_combout ))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[6][13]~q ),
	.datac(\storeregister[7][13]~q ),
	.datad(\Mux50~12_combout ),
	.cin(gnd),
	.combout(\Mux50~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~13 .lut_mask = 16'hF588;
defparam \Mux50~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N22
cycloneive_lcell_comb \Mux50~16 (
// Equation(s):
// \Mux50~16_combout  = (temp_imemload_output_19 & (((temp_imemload_output_18)))) # (!temp_imemload_output_19 & ((temp_imemload_output_18 & ((\Mux50~13_combout ))) # (!temp_imemload_output_18 & (\Mux50~15_combout ))))

	.dataa(\Mux50~15_combout ),
	.datab(temp_imemload_output_19),
	.datac(temp_imemload_output_18),
	.datad(\Mux50~13_combout ),
	.cin(gnd),
	.combout(\Mux50~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~16 .lut_mask = 16'hF2C2;
defparam \Mux50~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N8
cycloneive_lcell_comb \Mux50~17 (
// Equation(s):
// \Mux50~17_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & ((\storeregister[13][13]~q ))) # (!temp_imemload_output_16 & (\storeregister[12][13]~q ))))

	.dataa(\storeregister[12][13]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[13][13]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux50~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~17 .lut_mask = 16'hFC22;
defparam \Mux50~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N28
cycloneive_lcell_comb \Mux50~18 (
// Equation(s):
// \Mux50~18_combout  = (\Mux50~17_combout  & (((\storeregister[15][13]~q ) # (!temp_imemload_output_17)))) # (!\Mux50~17_combout  & (\storeregister[14][13]~q  & (temp_imemload_output_17)))

	.dataa(\storeregister[14][13]~q ),
	.datab(\Mux50~17_combout ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[15][13]~q ),
	.cin(gnd),
	.combout(\Mux50~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~18 .lut_mask = 16'hEC2C;
defparam \Mux50~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N4
cycloneive_lcell_comb \storeregister[27][11]~feeder (
// Equation(s):
// \storeregister[27][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux20),
	.datad(gnd),
	.cin(gnd),
	.combout(\storeregister[27][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[27][11]~feeder .lut_mask = 16'hF0F0;
defparam \storeregister[27][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N5
dffeas \storeregister[27][11] (
	.clk(!CLK),
	.d(\storeregister[27][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[27][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[27][11] .is_wysiwyg = "true";
defparam \storeregister[27][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N2
cycloneive_lcell_comb \Mux52~7 (
// Equation(s):
// \Mux52~7_combout  = (temp_imemload_output_18 & (((\storeregister[23][11]~q ) # (temp_imemload_output_19)))) # (!temp_imemload_output_18 & (\storeregister[19][11]~q  & ((!temp_imemload_output_19))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[19][11]~q ),
	.datac(\storeregister[23][11]~q ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux52~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~7 .lut_mask = 16'hAAE4;
defparam \Mux52~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N10
cycloneive_lcell_comb \Mux52~8 (
// Equation(s):
// \Mux52~8_combout  = (\Mux52~7_combout  & (((\storeregister[31][11]~q ) # (!temp_imemload_output_19)))) # (!\Mux52~7_combout  & (\storeregister[27][11]~q  & ((temp_imemload_output_19))))

	.dataa(\storeregister[27][11]~q ),
	.datab(\storeregister[31][11]~q ),
	.datac(\Mux52~7_combout ),
	.datad(temp_imemload_output_19),
	.cin(gnd),
	.combout(\Mux52~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~8 .lut_mask = 16'hCAF0;
defparam \Mux52~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N8
cycloneive_lcell_comb \Mux52~2 (
// Equation(s):
// \Mux52~2_combout  = (temp_imemload_output_19 & (((\storeregister[26][11]~q ) # (temp_imemload_output_18)))) # (!temp_imemload_output_19 & (\storeregister[18][11]~q  & ((!temp_imemload_output_18))))

	.dataa(temp_imemload_output_19),
	.datab(\storeregister[18][11]~q ),
	.datac(\storeregister[26][11]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux52~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~2 .lut_mask = 16'hAAE4;
defparam \Mux52~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N0
cycloneive_lcell_comb \Mux52~3 (
// Equation(s):
// \Mux52~3_combout  = (\Mux52~2_combout  & ((\storeregister[30][11]~q ) # ((!temp_imemload_output_18)))) # (!\Mux52~2_combout  & (((\storeregister[22][11]~q  & temp_imemload_output_18))))

	.dataa(\storeregister[30][11]~q ),
	.datab(\Mux52~2_combout ),
	.datac(\storeregister[22][11]~q ),
	.datad(temp_imemload_output_18),
	.cin(gnd),
	.combout(\Mux52~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~3 .lut_mask = 16'hB8CC;
defparam \Mux52~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N7
dffeas \storeregister[24][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[24][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[24][11] .is_wysiwyg = "true";
defparam \storeregister[24][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N6
cycloneive_lcell_comb \Mux52~4 (
// Equation(s):
// \Mux52~4_combout  = (temp_imemload_output_18 & (temp_imemload_output_19)) # (!temp_imemload_output_18 & ((temp_imemload_output_19 & (\storeregister[24][11]~q )) # (!temp_imemload_output_19 & ((\storeregister[16][11]~q )))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\storeregister[24][11]~q ),
	.datad(\storeregister[16][11]~q ),
	.cin(gnd),
	.combout(\Mux52~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~4 .lut_mask = 16'hD9C8;
defparam \Mux52~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N20
cycloneive_lcell_comb \storeregister[20][11]~feeder (
// Equation(s):
// \storeregister[20][11]~feeder_combout  = Mux20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux20),
	.cin(gnd),
	.combout(\storeregister[20][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \storeregister[20][11]~feeder .lut_mask = 16'hFF00;
defparam \storeregister[20][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N21
dffeas \storeregister[20][11] (
	.clk(!CLK),
	.d(\storeregister[20][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[20][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[20][11] .is_wysiwyg = "true";
defparam \storeregister[20][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N0
cycloneive_lcell_comb \Mux52~5 (
// Equation(s):
// \Mux52~5_combout  = (temp_imemload_output_18 & ((\Mux52~4_combout  & (\storeregister[28][11]~q )) # (!\Mux52~4_combout  & ((\storeregister[20][11]~q ))))) # (!temp_imemload_output_18 & (\Mux52~4_combout ))

	.dataa(temp_imemload_output_18),
	.datab(\Mux52~4_combout ),
	.datac(\storeregister[28][11]~q ),
	.datad(\storeregister[20][11]~q ),
	.cin(gnd),
	.combout(\Mux52~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~5 .lut_mask = 16'hE6C4;
defparam \Mux52~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N0
cycloneive_lcell_comb \Mux52~6 (
// Equation(s):
// \Mux52~6_combout  = (temp_imemload_output_16 & (((temp_imemload_output_17)))) # (!temp_imemload_output_16 & ((temp_imemload_output_17 & (\Mux52~3_combout )) # (!temp_imemload_output_17 & ((\Mux52~5_combout )))))

	.dataa(temp_imemload_output_16),
	.datab(\Mux52~3_combout ),
	.datac(temp_imemload_output_17),
	.datad(\Mux52~5_combout ),
	.cin(gnd),
	.combout(\Mux52~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~6 .lut_mask = 16'hE5E0;
defparam \Mux52~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N28
cycloneive_lcell_comb \Mux52~0 (
// Equation(s):
// \Mux52~0_combout  = (temp_imemload_output_18 & ((\storeregister[21][11]~q ) # ((temp_imemload_output_19)))) # (!temp_imemload_output_18 & (((!temp_imemload_output_19 & \storeregister[17][11]~q ))))

	.dataa(temp_imemload_output_18),
	.datab(\storeregister[21][11]~q ),
	.datac(temp_imemload_output_19),
	.datad(\storeregister[17][11]~q ),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~0 .lut_mask = 16'hADA8;
defparam \Mux52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N26
cycloneive_lcell_comb \Mux52~1 (
// Equation(s):
// \Mux52~1_combout  = (temp_imemload_output_19 & ((\Mux52~0_combout  & ((\storeregister[29][11]~q ))) # (!\Mux52~0_combout  & (\storeregister[25][11]~q )))) # (!temp_imemload_output_19 & (((\Mux52~0_combout ))))

	.dataa(\storeregister[25][11]~q ),
	.datab(\storeregister[29][11]~q ),
	.datac(temp_imemload_output_19),
	.datad(\Mux52~0_combout ),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~1 .lut_mask = 16'hCFA0;
defparam \Mux52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y42_N6
cycloneive_lcell_comb \Mux52~12 (
// Equation(s):
// \Mux52~12_combout  = (temp_imemload_output_17 & (((temp_imemload_output_16)))) # (!temp_imemload_output_17 & ((temp_imemload_output_16 & (\storeregister[5][11]~q )) # (!temp_imemload_output_16 & ((\storeregister[4][11]~q )))))

	.dataa(temp_imemload_output_17),
	.datab(\storeregister[5][11]~q ),
	.datac(\storeregister[4][11]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux52~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~12 .lut_mask = 16'hEE50;
defparam \Mux52~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N30
cycloneive_lcell_comb \Mux52~13 (
// Equation(s):
// \Mux52~13_combout  = (\Mux52~12_combout  & ((\storeregister[7][11]~q ) # ((!temp_imemload_output_17)))) # (!\Mux52~12_combout  & (((\storeregister[6][11]~q  & temp_imemload_output_17))))

	.dataa(\storeregister[7][11]~q ),
	.datab(\Mux52~12_combout ),
	.datac(\storeregister[6][11]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux52~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~13 .lut_mask = 16'hB8CC;
defparam \Mux52~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N14
cycloneive_lcell_comb \Mux52~15 (
// Equation(s):
// \Mux52~15_combout  = (\Mux52~14_combout ) # ((temp_imemload_output_17 & (\storeregister[2][11]~q  & !temp_imemload_output_16)))

	.dataa(\Mux52~14_combout ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[2][11]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux52~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~15 .lut_mask = 16'hAAEA;
defparam \Mux52~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N6
cycloneive_lcell_comb \Mux52~16 (
// Equation(s):
// \Mux52~16_combout  = (temp_imemload_output_18 & ((temp_imemload_output_19) # ((\Mux52~13_combout )))) # (!temp_imemload_output_18 & (!temp_imemload_output_19 & ((\Mux52~15_combout ))))

	.dataa(temp_imemload_output_18),
	.datab(temp_imemload_output_19),
	.datac(\Mux52~13_combout ),
	.datad(\Mux52~15_combout ),
	.cin(gnd),
	.combout(\Mux52~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~16 .lut_mask = 16'hB9A8;
defparam \Mux52~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N8
cycloneive_lcell_comb \Mux52~17 (
// Equation(s):
// \Mux52~17_combout  = (temp_imemload_output_16 & (((\storeregister[13][11]~q ) # (temp_imemload_output_17)))) # (!temp_imemload_output_16 & (\storeregister[12][11]~q  & ((!temp_imemload_output_17))))

	.dataa(\storeregister[12][11]~q ),
	.datab(temp_imemload_output_16),
	.datac(\storeregister[13][11]~q ),
	.datad(temp_imemload_output_17),
	.cin(gnd),
	.combout(\Mux52~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~17 .lut_mask = 16'hCCE2;
defparam \Mux52~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N24
cycloneive_lcell_comb \Mux52~18 (
// Equation(s):
// \Mux52~18_combout  = (\Mux52~17_combout  & (((\storeregister[15][11]~q ) # (!temp_imemload_output_17)))) # (!\Mux52~17_combout  & (\storeregister[14][11]~q  & (temp_imemload_output_17)))

	.dataa(\Mux52~17_combout ),
	.datab(\storeregister[14][11]~q ),
	.datac(temp_imemload_output_17),
	.datad(\storeregister[15][11]~q ),
	.cin(gnd),
	.combout(\Mux52~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~18 .lut_mask = 16'hEA4A;
defparam \Mux52~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y38_N17
dffeas \storeregister[10][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(Mux20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\storeregister[10][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \storeregister[10][11] .is_wysiwyg = "true";
defparam \storeregister[10][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N16
cycloneive_lcell_comb \Mux52~10 (
// Equation(s):
// \Mux52~10_combout  = (temp_imemload_output_17 & (((\storeregister[10][11]~q ) # (temp_imemload_output_16)))) # (!temp_imemload_output_17 & (\storeregister[8][11]~q  & ((!temp_imemload_output_16))))

	.dataa(\storeregister[8][11]~q ),
	.datab(temp_imemload_output_17),
	.datac(\storeregister[10][11]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux52~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~10 .lut_mask = 16'hCCE2;
defparam \Mux52~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N18
cycloneive_lcell_comb \Mux52~11 (
// Equation(s):
// \Mux52~11_combout  = (\Mux52~10_combout  & (((\storeregister[11][11]~q ) # (!temp_imemload_output_16)))) # (!\Mux52~10_combout  & (\storeregister[9][11]~q  & ((temp_imemload_output_16))))

	.dataa(\Mux52~10_combout ),
	.datab(\storeregister[9][11]~q ),
	.datac(\storeregister[11][11]~q ),
	.datad(temp_imemload_output_16),
	.cin(gnd),
	.combout(\Mux52~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~11 .lut_mask = 16'hE4AA;
defparam \Mux52~11 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module memory_control (
	temp_dmemWEN,
	temp_dmemREN,
	always1,
	ccifiwait_0,
	devpor,
	devclrn,
	devoe);
input 	temp_dmemWEN;
input 	temp_dmemREN;
input 	always1;
output 	ccifiwait_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X61_Y40_N4
cycloneive_lcell_comb \ccif.iwait[0]~0 (
// Equation(s):
// ccifiwait_0 = (temp_dmemREN1) # ((temp_dmemWEN1) # (!always1))

	.dataa(temp_dmemREN),
	.datab(always1),
	.datac(gnd),
	.datad(temp_dmemWEN),
	.cin(gnd),
	.combout(ccifiwait_0),
	.cout());
// synopsys translate_off
defparam \ccif.iwait[0]~0 .lut_mask = 16'hFFBB;
defparam \ccif.iwait[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module ram (
	is_in_use_reg,
	temp_dmemWEN,
	temp_dmemREN,
	ramaddr,
	ramaddr1,
	ramaddr2,
	ramaddr3,
	ramaddr4,
	ramaddr5,
	ramaddr6,
	ramaddr7,
	ramaddr8,
	ramaddr9,
	ramaddr10,
	ramaddr11,
	ramaddr12,
	ramaddr13,
	ramaddr14,
	ramaddr15,
	\ramif.ramaddr ,
	ramaddr16,
	ramaddr17,
	ramaddr18,
	ramaddr19,
	ramaddr20,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramWEN,
	ramstore,
	ramaddr21,
	ramaddr22,
	ramstore1,
	ramstore2,
	ramstore3,
	ramstore4,
	ramstore5,
	ramstore6,
	ramstore7,
	ramstore8,
	ramstore9,
	ramstore10,
	ramstore11,
	ramstore12,
	ramstore13,
	ramstore14,
	ramstore15,
	ramstore16,
	ramstore17,
	ramstore18,
	ramstore19,
	ramstore20,
	ramstore21,
	ramstore22,
	ramstore23,
	ramstore24,
	ramstore25,
	ramstore26,
	ramstore27,
	ramstore28,
	ramstore29,
	ramstore30,
	ramstore31,
	\ramif.ramREN ,
	ramaddr23,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	syifWEN,
	syiftbCTRL,
	syifREN,
	syifaddr_0,
	syifaddr_1,
	syifaddr_3,
	syifaddr_2,
	syifaddr_21,
	syifaddr_20,
	syifaddr_27,
	syifaddr_26,
	nRST,
	altera_internal_jtag1,
	nRST1,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	is_in_use_reg;
input 	temp_dmemWEN;
input 	temp_dmemREN;
input 	ramaddr;
input 	ramaddr1;
input 	ramaddr2;
input 	ramaddr3;
input 	ramaddr4;
input 	ramaddr5;
input 	ramaddr6;
input 	ramaddr7;
input 	ramaddr8;
input 	ramaddr9;
input 	ramaddr10;
input 	ramaddr11;
input 	ramaddr12;
input 	ramaddr13;
input 	ramaddr14;
input 	ramaddr15;
input 	[31:0] \ramif.ramaddr ;
input 	ramaddr16;
input 	ramaddr17;
input 	ramaddr18;
input 	ramaddr19;
input 	ramaddr20;
output 	always1;
output 	ramiframload_0;
output 	ramiframload_1;
output 	ramiframload_2;
output 	ramiframload_3;
output 	ramiframload_4;
output 	ramiframload_5;
output 	ramiframload_6;
output 	ramiframload_7;
output 	ramiframload_8;
output 	ramiframload_9;
output 	ramiframload_10;
output 	ramiframload_11;
output 	ramiframload_12;
output 	ramiframload_13;
output 	ramiframload_14;
output 	ramiframload_15;
output 	ramiframload_16;
output 	ramiframload_17;
output 	ramiframload_18;
output 	ramiframload_19;
output 	ramiframload_20;
output 	ramiframload_21;
output 	ramiframload_22;
output 	ramiframload_23;
output 	ramiframload_24;
output 	ramiframload_25;
output 	ramiframload_26;
output 	ramiframload_27;
output 	ramiframload_28;
output 	ramiframload_29;
output 	ramiframload_30;
output 	ramiframload_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramWEN;
input 	ramstore;
input 	ramaddr21;
input 	ramaddr22;
input 	ramstore1;
input 	ramstore2;
input 	ramstore3;
input 	ramstore4;
input 	ramstore5;
input 	ramstore6;
input 	ramstore7;
input 	ramstore8;
input 	ramstore9;
input 	ramstore10;
input 	ramstore11;
input 	ramstore12;
input 	ramstore13;
input 	ramstore14;
input 	ramstore15;
input 	ramstore16;
input 	ramstore17;
input 	ramstore18;
input 	ramstore19;
input 	ramstore20;
input 	ramstore21;
input 	ramstore22;
input 	ramstore23;
input 	ramstore24;
input 	ramstore25;
input 	ramstore26;
input 	ramstore27;
input 	ramstore28;
input 	ramstore29;
input 	ramstore30;
input 	ramstore31;
input 	\ramif.ramREN ;
input 	ramaddr23;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	syifWEN;
input 	syiftbCTRL;
input 	syifREN;
input 	syifaddr_0;
input 	syifaddr_1;
input 	syifaddr_3;
input 	syifaddr_2;
input 	syifaddr_21;
input 	syifaddr_20;
input 	syifaddr_27;
input 	syifaddr_26;
input 	nRST;
input 	altera_internal_jtag1;
input 	nRST1;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ;
wire \Equal2~0_combout ;
wire \Equal2~1_combout ;
wire \Equal2~2_combout ;
wire \Equal2~9_combout ;
wire \Equal2~10_combout ;
wire \Equal2~11_combout ;
wire \Equal2~12_combout ;
wire \Equal2~13_combout ;
wire \Equal2~17_combout ;
wire \Equal2~19_combout ;
wire \Equal2~22_combout ;
wire \Equal2~23_combout ;
wire \Equal2~24_combout ;
wire \always1~0_combout ;
wire \Equal2~4_combout ;
wire \Equal2~3_combout ;
wire \Equal2~5_combout ;
wire \Equal2~7_combout ;
wire \Equal2~6_combout ;
wire \Equal2~8_combout ;
wire \Equal2~26_combout ;
wire \Equal2~21_combout ;
wire \Equal2~25_combout ;
wire \Equal2~27_combout ;
wire \Equal2~16_combout ;
wire \Equal2~18_combout ;
wire \Equal2~14_combout ;
wire \Equal2~15_combout ;
wire \Equal2~20_combout ;
wire \Equal2~28_combout ;
wire \always0~3_combout ;
wire \always0~1_combout ;
wire \always0~0_combout ;
wire \always0~2_combout ;
wire \lcount~4_combout ;
wire \lcount~3_combout ;
wire \Add0~1_combout ;
wire \lcount~5_combout ;
wire \Add0~0_combout ;
wire \lcount~2_combout ;
wire \always1~1_combout ;
wire [3:0] lcount;
wire [1:0] en;
wire [31:0] addr;
wire [0:0] \altsyncram_component|auto_generated|altsyncram1|address_reg_a ;


altsyncram_1 altsyncram_component(
	.ram_block3a32(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.ram_block3a0(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.ram_block3a33(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.ram_block3a1(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.ram_block3a34(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.ram_block3a2(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.ram_block3a35(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.ram_block3a3(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.ram_block3a36(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.ram_block3a4(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.ram_block3a37(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.ram_block3a5(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.ram_block3a38(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.ram_block3a6(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.ram_block3a39(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.ram_block3a7(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.ram_block3a40(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.ram_block3a8(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.ram_block3a41(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.ram_block3a9(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.ram_block3a42(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.ram_block3a10(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.ram_block3a43(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.ram_block3a11(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.ram_block3a44(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.ram_block3a12(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.ram_block3a45(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.ram_block3a13(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.ram_block3a46(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.ram_block3a14(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.ram_block3a47(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.ram_block3a15(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.ram_block3a48(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.ram_block3a16(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.ram_block3a49(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.ram_block3a17(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.ram_block3a50(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.ram_block3a18(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.ram_block3a51(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.ram_block3a19(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.ram_block3a52(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.ram_block3a20(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.ram_block3a53(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.ram_block3a21(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.ram_block3a54(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.ram_block3a22(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.ram_block3a55(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.ram_block3a23(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.ram_block3a56(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.ram_block3a24(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.ram_block3a57(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.ram_block3a25(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.ram_block3a58(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.ram_block3a26(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.ram_block3a59(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.ram_block3a27(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.ram_block3a60(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.ram_block3a28(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.ram_block3a61(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.ram_block3a29(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.ram_block3a62(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.ram_block3a30(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.ram_block3a63(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.ram_block3a31(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.address_a({gnd,ramaddr15,ramaddr12,ramaddr13,ramaddr10,ramaddr11,ramaddr8,ramaddr9,ramaddr6,ramaddr7,ramaddr4,ramaddr5,ramaddr22,ramaddr21}),
	.ramaddr(ramaddr14),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.ramWEN(ramWEN),
	.data_a({ramstore31,ramstore30,ramstore29,ramstore28,ramstore27,ramstore26,ramstore25,ramstore24,ramstore23,ramstore22,ramstore21,ramstore20,ramstore19,ramstore18,ramstore17,ramstore16,ramstore15,ramstore14,ramstore13,ramstore12,ramstore11,ramstore10,ramstore9,ramstore8,ramstore7,ramstore6,
ramstore5,ramstore4,ramstore3,ramstore2,ramstore1,ramstore}),
	.ramaddr1(ramaddr23),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: FF_X63_Y43_N31
dffeas \addr[0] (
	.clk(!CLK),
	.d(\ramif.ramaddr [0]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[0] .is_wysiwyg = "true";
defparam \addr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N26
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = addr[0] $ (((\syif.tbCTRL~input_o  & (!\syif.addr[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((!\ramaddr~1_combout )))))

	.dataa(syiftbCTRL),
	.datab(syifaddr_0),
	.datac(addr[0]),
	.datad(ramaddr1),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'hD287;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y43_N1
dffeas \addr[1] (
	.clk(!CLK),
	.d(\ramif.ramaddr [1]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[1] .is_wysiwyg = "true";
defparam \addr[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N10
cycloneive_lcell_comb \Equal2~1 (
// Equation(s):
// \Equal2~1_combout  = addr[1] $ (((\syif.tbCTRL~input_o  & !\syif.addr[1]~input_o )))

	.dataa(syiftbCTRL),
	.datab(syifaddr_1),
	.datac(gnd),
	.datad(addr[1]),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~1 .lut_mask = 16'hDD22;
defparam \Equal2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N24
cycloneive_lcell_comb \Equal2~2 (
// Equation(s):
// \Equal2~2_combout  = (\Equal2~0_combout  & (\Equal2~1_combout  $ (((!\ramaddr~0_combout  & !\syif.tbCTRL~input_o )))))

	.dataa(ramaddr),
	.datab(syiftbCTRL),
	.datac(\Equal2~1_combout ),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~2 .lut_mask = 16'hE100;
defparam \Equal2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N5
dffeas \addr[4] (
	.clk(!CLK),
	.d(ramaddr5),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[4] .is_wysiwyg = "true";
defparam \addr[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N15
dffeas \addr[7] (
	.clk(!CLK),
	.d(ramaddr6),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[7] .is_wysiwyg = "true";
defparam \addr[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N27
dffeas \addr[8] (
	.clk(!CLK),
	.d(ramaddr9),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[8] .is_wysiwyg = "true";
defparam \addr[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N17
dffeas \addr[9] (
	.clk(!CLK),
	.d(ramaddr8),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[9] .is_wysiwyg = "true";
defparam \addr[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N6
cycloneive_lcell_comb \Equal2~9 (
// Equation(s):
// \Equal2~9_combout  = (addr[9] & (\ramaddr~13_combout  & (addr[8] $ (!\ramaddr~15_combout )))) # (!addr[9] & (!\ramaddr~13_combout  & (addr[8] $ (!\ramaddr~15_combout ))))

	.dataa(addr[9]),
	.datab(addr[8]),
	.datac(ramaddr9),
	.datad(ramaddr8),
	.cin(gnd),
	.combout(\Equal2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~9 .lut_mask = 16'h8241;
defparam \Equal2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y43_N25
dffeas \addr[10] (
	.clk(!CLK),
	.d(ramaddr11),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[10] .is_wysiwyg = "true";
defparam \addr[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y43_N15
dffeas \addr[11] (
	.clk(!CLK),
	.d(ramaddr10),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[11] .is_wysiwyg = "true";
defparam \addr[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N4
cycloneive_lcell_comb \Equal2~10 (
// Equation(s):
// \Equal2~10_combout  = (addr[10] & (\ramaddr~19_combout  & (addr[11] $ (!\ramaddr~17_combout )))) # (!addr[10] & (!\ramaddr~19_combout  & (addr[11] $ (!\ramaddr~17_combout ))))

	.dataa(addr[10]),
	.datab(addr[11]),
	.datac(ramaddr10),
	.datad(ramaddr11),
	.cin(gnd),
	.combout(\Equal2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~10 .lut_mask = 16'h8241;
defparam \Equal2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y43_N23
dffeas \addr[12] (
	.clk(!CLK),
	.d(ramaddr13),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[12] .is_wysiwyg = "true";
defparam \addr[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y43_N9
dffeas \addr[13] (
	.clk(!CLK),
	.d(ramaddr12),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[13] .is_wysiwyg = "true";
defparam \addr[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N0
cycloneive_lcell_comb \Equal2~11 (
// Equation(s):
// \Equal2~11_combout  = (addr[13] & (\ramaddr~21_combout  & (addr[12] $ (!\ramaddr~23_combout )))) # (!addr[13] & (!\ramaddr~21_combout  & (addr[12] $ (!\ramaddr~23_combout ))))

	.dataa(addr[13]),
	.datab(addr[12]),
	.datac(ramaddr13),
	.datad(ramaddr12),
	.cin(gnd),
	.combout(\Equal2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~11 .lut_mask = 16'h8241;
defparam \Equal2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y43_N23
dffeas \addr[14] (
	.clk(!CLK),
	.d(ramaddr15),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[14] .is_wysiwyg = "true";
defparam \addr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N21
dffeas \addr[15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(ramaddr23),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[15] .is_wysiwyg = "true";
defparam \addr[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N26
cycloneive_lcell_comb \Equal2~12 (
// Equation(s):
// \Equal2~12_combout  = (addr[14] & (\ramaddr~27_combout  & (addr[15] $ (\ramaddr~25_combout )))) # (!addr[14] & (!\ramaddr~27_combout  & (addr[15] $ (\ramaddr~25_combout ))))

	.dataa(addr[14]),
	.datab(addr[15]),
	.datac(ramaddr15),
	.datad(ramaddr14),
	.cin(gnd),
	.combout(\Equal2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~12 .lut_mask = 16'h2184;
defparam \Equal2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N12
cycloneive_lcell_comb \Equal2~13 (
// Equation(s):
// \Equal2~13_combout  = (\Equal2~9_combout  & (\Equal2~11_combout  & (\Equal2~12_combout  & \Equal2~10_combout )))

	.dataa(\Equal2~9_combout ),
	.datab(\Equal2~11_combout ),
	.datac(\Equal2~12_combout ),
	.datad(\Equal2~10_combout ),
	.cin(gnd),
	.combout(\Equal2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~13 .lut_mask = 16'h8000;
defparam \Equal2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y43_N9
dffeas \addr[17] (
	.clk(!CLK),
	.d(\ramif.ramaddr [17]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[17]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[17] .is_wysiwyg = "true";
defparam \addr[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y43_N21
dffeas \addr[19] (
	.clk(!CLK),
	.d(\ramif.ramaddr [19]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[19] .is_wysiwyg = "true";
defparam \addr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y43_N17
dffeas \addr[20] (
	.clk(!CLK),
	.d(\ramif.ramaddr [20]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[20] .is_wysiwyg = "true";
defparam \addr[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N14
cycloneive_lcell_comb \Equal2~17 (
// Equation(s):
// \Equal2~17_combout  = addr[20] $ (((\syif.tbCTRL~input_o  & !\syif.addr[20]~input_o )))

	.dataa(syiftbCTRL),
	.datab(syifaddr_20),
	.datac(gnd),
	.datad(addr[20]),
	.cin(gnd),
	.combout(\Equal2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~17 .lut_mask = 16'hDD22;
defparam \Equal2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N9
dffeas \addr[22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(ramaddr18),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[22] .is_wysiwyg = "true";
defparam \addr[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N15
dffeas \addr[23] (
	.clk(!CLK),
	.d(\ramif.ramaddr [23]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[23] .is_wysiwyg = "true";
defparam \addr[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N6
cycloneive_lcell_comb \Equal2~19 (
// Equation(s):
// \Equal2~19_combout  = (addr[23] & (\ramaddr~39_combout  & (addr[22] $ (!\ramaddr~41_combout )))) # (!addr[23] & (!\ramaddr~39_combout  & (addr[22] $ (!\ramaddr~41_combout ))))

	.dataa(addr[23]),
	.datab(addr[22]),
	.datac(\ramif.ramaddr [23]),
	.datad(ramaddr18),
	.cin(gnd),
	.combout(\Equal2~19_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~19 .lut_mask = 16'h8421;
defparam \Equal2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y43_N25
dffeas \addr[24] (
	.clk(!CLK),
	.d(\ramif.ramaddr [24]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[24] .is_wysiwyg = "true";
defparam \addr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y43_N31
dffeas \addr[27] (
	.clk(!CLK),
	.d(\ramif.ramaddr [27]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[27]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[27] .is_wysiwyg = "true";
defparam \addr[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N10
cycloneive_lcell_comb \Equal2~22 (
// Equation(s):
// \Equal2~22_combout  = addr[27] $ (((\syif.tbCTRL~input_o  & (!\syif.addr[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((!\ramaddr~47_combout )))))

	.dataa(syiftbCTRL),
	.datab(addr[27]),
	.datac(syifaddr_27),
	.datad(ramaddr20),
	.cin(gnd),
	.combout(\Equal2~22_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~22 .lut_mask = 16'hC693;
defparam \Equal2~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y43_N17
dffeas \addr[26] (
	.clk(!CLK),
	.d(\ramif.ramaddr [26]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[26]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[26] .is_wysiwyg = "true";
defparam \addr[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N4
cycloneive_lcell_comb \Equal2~23 (
// Equation(s):
// \Equal2~23_combout  = addr[26] $ (((!\syif.addr[26]~input_o  & \syif.tbCTRL~input_o )))

	.dataa(syifaddr_26),
	.datab(syiftbCTRL),
	.datac(gnd),
	.datad(addr[26]),
	.cin(gnd),
	.combout(\Equal2~23_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~23 .lut_mask = 16'hBB44;
defparam \Equal2~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N22
cycloneive_lcell_comb \Equal2~24 (
// Equation(s):
// \Equal2~24_combout  = (\Equal2~22_combout  & (\Equal2~23_combout  $ (((!\syif.tbCTRL~input_o  & !\ramaddr~46_combout )))))

	.dataa(syiftbCTRL),
	.datab(\Equal2~23_combout ),
	.datac(ramaddr19),
	.datad(\Equal2~22_combout ),
	.cin(gnd),
	.combout(\Equal2~24_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~24 .lut_mask = 16'hC900;
defparam \Equal2~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y43_N29
dffeas \addr[30] (
	.clk(!CLK),
	.d(\ramif.ramaddr [30]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[30]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[30] .is_wysiwyg = "true";
defparam \addr[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N7
dffeas \en[1] (
	.clk(!CLK),
	.d(\ramif.ramREN ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[1]),
	.prn(vcc));
// synopsys translate_off
defparam \en[1] .is_wysiwyg = "true";
defparam \en[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N30
cycloneive_lcell_comb \always1~2 (
// Equation(s):
// always1 = ((!\always1~0_combout  & (\always1~1_combout  & \Equal2~28_combout ))) # (!\nRST~input_o )

	.dataa(\always1~0_combout ),
	.datab(\always1~1_combout ),
	.datac(nRST),
	.datad(\Equal2~28_combout ),
	.cin(gnd),
	.combout(always1),
	.cout());
// synopsys translate_off
defparam \always1~2 .lut_mask = 16'h4F0F;
defparam \always1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N16
cycloneive_lcell_comb \ramif.ramload[0]~0 (
// Equation(s):
// ramiframload_0 = ((address_reg_a_0 & ((ram_block3a321))) # (!address_reg_a_0 & (ram_block3a01))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.cin(gnd),
	.combout(ramiframload_0),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~0 .lut_mask = 16'hFD5D;
defparam \ramif.ramload[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y40_N20
cycloneive_lcell_comb \ramif.ramload[1]~1 (
// Equation(s):
// ramiframload_1 = (always1 & ((address_reg_a_0 & ((ram_block3a331))) # (!address_reg_a_0 & (ram_block3a110))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.cin(gnd),
	.combout(ramiframload_1),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[1]~1 .lut_mask = 16'hA808;
defparam \ramif.ramload[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N16
cycloneive_lcell_comb \ramif.ramload[2]~2 (
// Equation(s):
// ramiframload_2 = (always1 & ((address_reg_a_0 & (ram_block3a341)) # (!address_reg_a_0 & ((ram_block3a210)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_2),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[2]~2 .lut_mask = 16'hA0C0;
defparam \ramif.ramload[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y40_N22
cycloneive_lcell_comb \ramif.ramload[3]~3 (
// Equation(s):
// ramiframload_3 = (always1 & ((address_reg_a_0 & (ram_block3a351)) # (!address_reg_a_0 & ((ram_block3a310)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.cin(gnd),
	.combout(ramiframload_3),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[3]~3 .lut_mask = 16'h8A80;
defparam \ramif.ramload[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N24
cycloneive_lcell_comb \ramif.ramload[4]~4 (
// Equation(s):
// ramiframload_4 = ((address_reg_a_0 & (ram_block3a361)) # (!address_reg_a_0 & ((ram_block3a410)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.cin(gnd),
	.combout(ramiframload_4),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[4]~4 .lut_mask = 16'hDF8F;
defparam \ramif.ramload[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N26
cycloneive_lcell_comb \ramif.ramload[5]~5 (
// Equation(s):
// ramiframload_5 = (always1 & ((address_reg_a_0 & ((ram_block3a371))) # (!address_reg_a_0 & (ram_block3a510))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_5),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[5]~5 .lut_mask = 16'hC0A0;
defparam \ramif.ramload[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N26
cycloneive_lcell_comb \ramif.ramload[6]~6 (
// Equation(s):
// ramiframload_6 = ((address_reg_a_0 & (ram_block3a381)) # (!address_reg_a_0 & ((ram_block3a64)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_6),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[6]~6 .lut_mask = 16'hACFF;
defparam \ramif.ramload[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N16
cycloneive_lcell_comb \ramif.ramload[7]~7 (
// Equation(s):
// ramiframload_7 = ((address_reg_a_0 & (ram_block3a391)) # (!address_reg_a_0 & ((ram_block3a71)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.cin(gnd),
	.combout(ramiframload_7),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[7]~7 .lut_mask = 16'hBF8F;
defparam \ramif.ramload[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y40_N0
cycloneive_lcell_comb \ramif.ramload[8]~8 (
// Equation(s):
// ramiframload_8 = (always1 & ((address_reg_a_0 & ((ram_block3a401))) # (!address_reg_a_0 & (ram_block3a81))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.cin(gnd),
	.combout(ramiframload_8),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[8]~8 .lut_mask = 16'hE020;
defparam \ramif.ramload[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y40_N6
cycloneive_lcell_comb \ramif.ramload[9]~9 (
// Equation(s):
// ramiframload_9 = ((address_reg_a_0 & (ram_block3a412)) # (!address_reg_a_0 & ((ram_block3a91)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.cin(gnd),
	.combout(ramiframload_9),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[9]~9 .lut_mask = 16'hDFD5;
defparam \ramif.ramload[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y40_N12
cycloneive_lcell_comb \ramif.ramload[10]~10 (
// Equation(s):
// ramiframload_10 = (always1 & ((address_reg_a_0 & (ram_block3a421)) # (!address_reg_a_0 & ((ram_block3a101)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.cin(gnd),
	.combout(ramiframload_10),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[10]~10 .lut_mask = 16'hB080;
defparam \ramif.ramload[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N18
cycloneive_lcell_comb \ramif.ramload[11]~11 (
// Equation(s):
// ramiframload_11 = ((address_reg_a_0 & ((ram_block3a431))) # (!address_reg_a_0 & (ram_block3a112))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_11),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[11]~11 .lut_mask = 16'hF5DD;
defparam \ramif.ramload[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y40_N26
cycloneive_lcell_comb \ramif.ramload[12]~12 (
// Equation(s):
// ramiframload_12 = ((address_reg_a_0 & ((ram_block3a441))) # (!address_reg_a_0 & (ram_block3a121))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.cin(gnd),
	.combout(ramiframload_12),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[12]~12 .lut_mask = 16'hFD5D;
defparam \ramif.ramload[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y40_N4
cycloneive_lcell_comb \ramif.ramload[13]~13 (
// Equation(s):
// ramiframload_13 = ((address_reg_a_0 & (ram_block3a451)) # (!address_reg_a_0 & ((ram_block3a131)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.cin(gnd),
	.combout(ramiframload_13),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[13]~13 .lut_mask = 16'hDFD5;
defparam \ramif.ramload[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y40_N30
cycloneive_lcell_comb \ramif.ramload[14]~14 (
// Equation(s):
// ramiframload_14 = (always1 & ((address_reg_a_0 & (ram_block3a461)) # (!address_reg_a_0 & ((ram_block3a141)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.cin(gnd),
	.combout(ramiframload_14),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[14]~14 .lut_mask = 16'hB080;
defparam \ramif.ramload[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N12
cycloneive_lcell_comb \ramif.ramload[15]~15 (
// Equation(s):
// ramiframload_15 = ((address_reg_a_0 & (ram_block3a471)) # (!address_reg_a_0 & ((ram_block3a151)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_15),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[15]~15 .lut_mask = 16'hD8FF;
defparam \ramif.ramload[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N12
cycloneive_lcell_comb \ramif.ramload[16]~16 (
// Equation(s):
// ramiframload_16 = ((address_reg_a_0 & (ram_block3a481)) # (!address_reg_a_0 & ((ram_block3a161)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_16),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[16]~16 .lut_mask = 16'hD8FF;
defparam \ramif.ramload[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N2
cycloneive_lcell_comb \ramif.ramload[17]~17 (
// Equation(s):
// ramiframload_17 = (always1 & ((address_reg_a_0 & (ram_block3a491)) # (!address_reg_a_0 & ((ram_block3a171)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_17),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[17]~17 .lut_mask = 16'hD800;
defparam \ramif.ramload[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N8
cycloneive_lcell_comb \ramif.ramload[18]~18 (
// Equation(s):
// ramiframload_18 = (always1 & ((address_reg_a_0 & ((ram_block3a501))) # (!address_reg_a_0 & (ram_block3a181))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_18),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[18]~18 .lut_mask = 16'hE400;
defparam \ramif.ramload[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N14
cycloneive_lcell_comb \ramif.ramload[19]~19 (
// Equation(s):
// ramiframload_19 = (always1 & ((address_reg_a_0 & (ram_block3a512)) # (!address_reg_a_0 & ((ram_block3a191)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_19),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[19]~19 .lut_mask = 16'hAC00;
defparam \ramif.ramload[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N24
cycloneive_lcell_comb \ramif.ramload[20]~20 (
// Equation(s):
// ramiframload_20 = ((address_reg_a_0 & (ram_block3a521)) # (!address_reg_a_0 & ((ram_block3a201)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.cin(gnd),
	.combout(ramiframload_20),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[20]~20 .lut_mask = 16'hBF8F;
defparam \ramif.ramload[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N20
cycloneive_lcell_comb \ramif.ramload[21]~21 (
// Equation(s):
// ramiframload_21 = (always1 & ((address_reg_a_0 & ((ram_block3a531))) # (!address_reg_a_0 & (ram_block3a212))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_21),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[21]~21 .lut_mask = 16'hCA00;
defparam \ramif.ramload[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N6
cycloneive_lcell_comb \ramif.ramload[22]~22 (
// Equation(s):
// ramiframload_22 = ((address_reg_a_0 & (ram_block3a541)) # (!address_reg_a_0 & ((ram_block3a221)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_22),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[22]~22 .lut_mask = 16'hACFF;
defparam \ramif.ramload[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N24
cycloneive_lcell_comb \ramif.ramload[23]~23 (
// Equation(s):
// ramiframload_23 = ((address_reg_a_0 & ((ram_block3a551))) # (!address_reg_a_0 & (ram_block3a231))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_23),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[23]~23 .lut_mask = 16'hCAFF;
defparam \ramif.ramload[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N18
cycloneive_lcell_comb \ramif.ramload[24]~24 (
// Equation(s):
// ramiframload_24 = (always1 & ((address_reg_a_0 & ((ram_block3a561))) # (!address_reg_a_0 & (ram_block3a241))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_24),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[24]~24 .lut_mask = 16'hCA00;
defparam \ramif.ramload[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N28
cycloneive_lcell_comb \ramif.ramload[25]~25 (
// Equation(s):
// ramiframload_25 = ((address_reg_a_0 & ((ram_block3a571))) # (!address_reg_a_0 & (ram_block3a251))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_25),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[25]~25 .lut_mask = 16'hCAFF;
defparam \ramif.ramload[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N30
cycloneive_lcell_comb \ramif.ramload[26]~26 (
// Equation(s):
// ramiframload_26 = (always1 & ((address_reg_a_0 & (ram_block3a581)) # (!address_reg_a_0 & ((ram_block3a261)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_26),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[26]~26 .lut_mask = 16'hD800;
defparam \ramif.ramload[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N16
cycloneive_lcell_comb \ramif.ramload[27]~27 (
// Equation(s):
// ramiframload_27 = ((address_reg_a_0 & ((ram_block3a591))) # (!address_reg_a_0 & (ram_block3a271))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_27),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[27]~27 .lut_mask = 16'hE4FF;
defparam \ramif.ramload[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N4
cycloneive_lcell_comb \ramif.ramload[28]~28 (
// Equation(s):
// ramiframload_28 = ((address_reg_a_0 & ((ram_block3a601))) # (!address_reg_a_0 & (ram_block3a281))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.cin(gnd),
	.combout(ramiframload_28),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[28]~28 .lut_mask = 16'hEF4F;
defparam \ramif.ramload[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N16
cycloneive_lcell_comb \ramif.ramload[29]~29 (
// Equation(s):
// ramiframload_29 = ((address_reg_a_0 & (ram_block3a611)) # (!address_reg_a_0 & ((ram_block3a291)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_29),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[29]~29 .lut_mask = 16'hD8FF;
defparam \ramif.ramload[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N18
cycloneive_lcell_comb \ramif.ramload[30]~30 (
// Equation(s):
// ramiframload_30 = (always1 & ((address_reg_a_0 & (ram_block3a621)) # (!address_reg_a_0 & ((ram_block3a301)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.cin(gnd),
	.combout(ramiframload_30),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[30]~30 .lut_mask = 16'hA280;
defparam \ramif.ramload[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N28
cycloneive_lcell_comb \ramif.ramload[31]~31 (
// Equation(s):
// ramiframload_31 = ((address_reg_a_0 & (ram_block3a631)) # (!address_reg_a_0 & ((ram_block3a312)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.cin(gnd),
	.combout(ramiframload_31),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[31]~31 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N12
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// \always1~0_combout  = (!\syif.WEN~input_o  & (\syif.tbCTRL~input_o  & !\syif.REN~input_o ))

	.dataa(gnd),
	.datab(syifWEN),
	.datac(syiftbCTRL),
	.datad(syifREN),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'h0030;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N19
dffeas \addr[2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(ramaddr21),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[2] .is_wysiwyg = "true";
defparam \addr[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N18
cycloneive_lcell_comb \Equal2~4 (
// Equation(s):
// \Equal2~4_combout  = addr[2] $ (((\syif.tbCTRL~input_o  & !\syif.addr[2]~input_o )))

	.dataa(syiftbCTRL),
	.datab(gnd),
	.datac(addr[2]),
	.datad(syifaddr_2),
	.cin(gnd),
	.combout(\Equal2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~4 .lut_mask = 16'hF05A;
defparam \Equal2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N31
dffeas \addr[3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(ramaddr22),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[3] .is_wysiwyg = "true";
defparam \addr[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N30
cycloneive_lcell_comb \Equal2~3 (
// Equation(s):
// \Equal2~3_combout  = addr[3] $ (((\syif.tbCTRL~input_o  & (!\syif.addr[3]~input_o )) # (!\syif.tbCTRL~input_o  & ((!\ramaddr~3_combout )))))

	.dataa(syiftbCTRL),
	.datab(syifaddr_3),
	.datac(addr[3]),
	.datad(ramaddr3),
	.cin(gnd),
	.combout(\Equal2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~3 .lut_mask = 16'hD287;
defparam \Equal2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N24
cycloneive_lcell_comb \Equal2~5 (
// Equation(s):
// \Equal2~5_combout  = (\Equal2~3_combout  & (\Equal2~4_combout  $ (((!\syif.tbCTRL~input_o  & !\ramaddr~2_combout )))))

	.dataa(syiftbCTRL),
	.datab(\Equal2~4_combout ),
	.datac(\Equal2~3_combout ),
	.datad(ramaddr2),
	.cin(gnd),
	.combout(\Equal2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~5 .lut_mask = 16'hC090;
defparam \Equal2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y43_N13
dffeas \addr[6] (
	.clk(!CLK),
	.d(ramaddr7),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[6] .is_wysiwyg = "true";
defparam \addr[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N4
cycloneive_lcell_comb \Equal2~7 (
// Equation(s):
// \Equal2~7_combout  = (addr[7] & (\ramaddr~9_combout  & (addr[6] $ (!\ramaddr~11_combout )))) # (!addr[7] & (!\ramaddr~9_combout  & (addr[6] $ (!\ramaddr~11_combout ))))

	.dataa(addr[7]),
	.datab(addr[6]),
	.datac(ramaddr6),
	.datad(ramaddr7),
	.cin(gnd),
	.combout(\Equal2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~7 .lut_mask = 16'h8421;
defparam \Equal2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N19
dffeas \addr[5] (
	.clk(!CLK),
	.d(ramaddr4),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[5] .is_wysiwyg = "true";
defparam \addr[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N0
cycloneive_lcell_comb \Equal2~6 (
// Equation(s):
// \Equal2~6_combout  = (addr[4] & (\ramaddr~7_combout  & (addr[5] $ (!\ramaddr~5_combout )))) # (!addr[4] & (!\ramaddr~7_combout  & (addr[5] $ (!\ramaddr~5_combout ))))

	.dataa(addr[4]),
	.datab(addr[5]),
	.datac(ramaddr5),
	.datad(ramaddr4),
	.cin(gnd),
	.combout(\Equal2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~6 .lut_mask = 16'h8421;
defparam \Equal2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N2
cycloneive_lcell_comb \Equal2~8 (
// Equation(s):
// \Equal2~8_combout  = (\Equal2~2_combout  & (\Equal2~5_combout  & (\Equal2~7_combout  & \Equal2~6_combout )))

	.dataa(\Equal2~2_combout ),
	.datab(\Equal2~5_combout ),
	.datac(\Equal2~7_combout ),
	.datad(\Equal2~6_combout ),
	.cin(gnd),
	.combout(\Equal2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~8 .lut_mask = 16'h8000;
defparam \Equal2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y43_N31
dffeas \addr[31] (
	.clk(!CLK),
	.d(\ramif.ramaddr [31]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[31]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[31] .is_wysiwyg = "true";
defparam \addr[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N24
cycloneive_lcell_comb \Equal2~26 (
// Equation(s):
// \Equal2~26_combout  = (addr[30] & (\ramaddr~55_combout  & (addr[31] $ (!\ramaddr~53_combout )))) # (!addr[30] & (!\ramaddr~55_combout  & (addr[31] $ (!\ramaddr~53_combout ))))

	.dataa(addr[30]),
	.datab(addr[31]),
	.datac(\ramif.ramaddr [31]),
	.datad(\ramif.ramaddr [30]),
	.cin(gnd),
	.combout(\Equal2~26_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~26 .lut_mask = 16'h8241;
defparam \Equal2~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y43_N19
dffeas \addr[25] (
	.clk(!CLK),
	.d(\ramif.ramaddr [25]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[25] .is_wysiwyg = "true";
defparam \addr[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N14
cycloneive_lcell_comb \Equal2~21 (
// Equation(s):
// \Equal2~21_combout  = (addr[24] & (\ramaddr~45_combout  & (\ramaddr~43_combout  $ (!addr[25])))) # (!addr[24] & (!\ramaddr~45_combout  & (\ramaddr~43_combout  $ (!addr[25]))))

	.dataa(addr[24]),
	.datab(\ramif.ramaddr [25]),
	.datac(addr[25]),
	.datad(\ramif.ramaddr [24]),
	.cin(gnd),
	.combout(\Equal2~21_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~21 .lut_mask = 16'h8241;
defparam \Equal2~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y43_N13
dffeas \addr[28] (
	.clk(!CLK),
	.d(\ramif.ramaddr [28]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[28]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[28] .is_wysiwyg = "true";
defparam \addr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y43_N7
dffeas \addr[29] (
	.clk(!CLK),
	.d(\ramif.ramaddr [29]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[29]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[29] .is_wysiwyg = "true";
defparam \addr[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N26
cycloneive_lcell_comb \Equal2~25 (
// Equation(s):
// \Equal2~25_combout  = (\ramaddr~51_combout  & (addr[28] & (addr[29] $ (!\ramaddr~49_combout )))) # (!\ramaddr~51_combout  & (!addr[28] & (addr[29] $ (!\ramaddr~49_combout ))))

	.dataa(\ramif.ramaddr [28]),
	.datab(addr[28]),
	.datac(addr[29]),
	.datad(\ramif.ramaddr [29]),
	.cin(gnd),
	.combout(\Equal2~25_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~25 .lut_mask = 16'h9009;
defparam \Equal2~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N26
cycloneive_lcell_comb \Equal2~27 (
// Equation(s):
// \Equal2~27_combout  = (\Equal2~24_combout  & (\Equal2~26_combout  & (\Equal2~21_combout  & \Equal2~25_combout )))

	.dataa(\Equal2~24_combout ),
	.datab(\Equal2~26_combout ),
	.datac(\Equal2~21_combout ),
	.datad(\Equal2~25_combout ),
	.cin(gnd),
	.combout(\Equal2~27_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~27 .lut_mask = 16'h8000;
defparam \Equal2~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y43_N5
dffeas \addr[21] (
	.clk(!CLK),
	.d(\ramif.ramaddr [21]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[21] .is_wysiwyg = "true";
defparam \addr[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N10
cycloneive_lcell_comb \Equal2~16 (
// Equation(s):
// \Equal2~16_combout  = addr[21] $ (((\syif.tbCTRL~input_o  & (!\syif.addr[21]~input_o )) # (!\syif.tbCTRL~input_o  & ((!\ramaddr~37_combout )))))

	.dataa(syiftbCTRL),
	.datab(syifaddr_21),
	.datac(addr[21]),
	.datad(ramaddr17),
	.cin(gnd),
	.combout(\Equal2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~16 .lut_mask = 16'hD287;
defparam \Equal2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N6
cycloneive_lcell_comb \Equal2~18 (
// Equation(s):
// \Equal2~18_combout  = (\Equal2~16_combout  & (\Equal2~17_combout  $ (((!\ramaddr~36_combout  & !\syif.tbCTRL~input_o )))))

	.dataa(\Equal2~17_combout ),
	.datab(ramaddr16),
	.datac(syiftbCTRL),
	.datad(\Equal2~16_combout ),
	.cin(gnd),
	.combout(\Equal2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~18 .lut_mask = 16'hA900;
defparam \Equal2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y43_N11
dffeas \addr[16] (
	.clk(!CLK),
	.d(\ramif.ramaddr [16]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[16]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[16] .is_wysiwyg = "true";
defparam \addr[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N28
cycloneive_lcell_comb \Equal2~14 (
// Equation(s):
// \Equal2~14_combout  = (addr[17] & (\ramaddr~29_combout  & (addr[16] $ (!\ramaddr~31_combout )))) # (!addr[17] & (!\ramaddr~29_combout  & (addr[16] $ (!\ramaddr~31_combout ))))

	.dataa(addr[17]),
	.datab(addr[16]),
	.datac(\ramif.ramaddr [17]),
	.datad(\ramif.ramaddr [16]),
	.cin(gnd),
	.combout(\Equal2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~14 .lut_mask = 16'h8421;
defparam \Equal2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y43_N31
dffeas \addr[18] (
	.clk(!CLK),
	.d(\ramif.ramaddr [18]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[18] .is_wysiwyg = "true";
defparam \addr[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N22
cycloneive_lcell_comb \Equal2~15 (
// Equation(s):
// \Equal2~15_combout  = (addr[19] & (\ramaddr~33_combout  & (addr[18] $ (!\ramaddr~35_combout )))) # (!addr[19] & (!\ramaddr~33_combout  & (addr[18] $ (!\ramaddr~35_combout ))))

	.dataa(addr[19]),
	.datab(addr[18]),
	.datac(\ramif.ramaddr [18]),
	.datad(\ramif.ramaddr [19]),
	.cin(gnd),
	.combout(\Equal2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~15 .lut_mask = 16'h8241;
defparam \Equal2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N24
cycloneive_lcell_comb \Equal2~20 (
// Equation(s):
// \Equal2~20_combout  = (\Equal2~19_combout  & (\Equal2~18_combout  & (\Equal2~14_combout  & \Equal2~15_combout )))

	.dataa(\Equal2~19_combout ),
	.datab(\Equal2~18_combout ),
	.datac(\Equal2~14_combout ),
	.datad(\Equal2~15_combout ),
	.cin(gnd),
	.combout(\Equal2~20_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~20 .lut_mask = 16'h8000;
defparam \Equal2~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N28
cycloneive_lcell_comb \Equal2~28 (
// Equation(s):
// \Equal2~28_combout  = (\Equal2~13_combout  & (\Equal2~8_combout  & (\Equal2~27_combout  & \Equal2~20_combout )))

	.dataa(\Equal2~13_combout ),
	.datab(\Equal2~8_combout ),
	.datac(\Equal2~27_combout ),
	.datad(\Equal2~20_combout ),
	.cin(gnd),
	.combout(\Equal2~28_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~28 .lut_mask = 16'h8000;
defparam \Equal2~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N14
cycloneive_lcell_comb \always0~3 (
// Equation(s):
// \always0~3_combout  = (\always0~2_combout ) # ((\always1~0_combout ) # (!\Equal2~28_combout ))

	.dataa(gnd),
	.datab(\always0~2_combout ),
	.datac(\always1~0_combout ),
	.datad(\Equal2~28_combout ),
	.cin(gnd),
	.combout(\always0~3_combout ),
	.cout());
// synopsys translate_off
defparam \always0~3 .lut_mask = 16'hFCFF;
defparam \always0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N23
dffeas \en[0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(ramWEN),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[0]),
	.prn(vcc));
// synopsys translate_off
defparam \en[0] .is_wysiwyg = "true";
defparam \en[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N24
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = en[0] $ (((\syif.WEN~input_o  & \syif.tbCTRL~input_o )))

	.dataa(gnd),
	.datab(syifWEN),
	.datac(syiftbCTRL),
	.datad(en[0]),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'h3FC0;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N2
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (\syif.tbCTRL~input_o  & (((\syif.REN~input_o )))) # (!\syif.tbCTRL~input_o  & (!temp_dmemREN1 & ((temp_dmemWEN1))))

	.dataa(temp_dmemREN),
	.datab(syifREN),
	.datac(temp_dmemWEN),
	.datad(syiftbCTRL),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'hCC50;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N10
cycloneive_lcell_comb \always0~2 (
// Equation(s):
// \always0~2_combout  = (en[1] & ((\always0~1_combout ) # (\syif.tbCTRL~input_o  $ (\always0~0_combout )))) # (!en[1] & ((\always0~1_combout  & ((\syif.tbCTRL~input_o ) # (!\always0~0_combout ))) # (!\always0~1_combout  & ((\always0~0_combout ) # 
// (!\syif.tbCTRL~input_o )))))

	.dataa(en[1]),
	.datab(\always0~1_combout ),
	.datac(syiftbCTRL),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
// synopsys translate_off
defparam \always0~2 .lut_mask = 16'hDBED;
defparam \always0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N10
cycloneive_lcell_comb \lcount~4 (
// Equation(s):
// \lcount~4_combout  = (\always1~0_combout ) # ((\always0~2_combout ) # ((!\Equal2~28_combout ) # (!lcount[0])))

	.dataa(\always1~0_combout ),
	.datab(\always0~2_combout ),
	.datac(lcount[0]),
	.datad(\Equal2~28_combout ),
	.cin(gnd),
	.combout(\lcount~4_combout ),
	.cout());
// synopsys translate_off
defparam \lcount~4 .lut_mask = 16'hEFFF;
defparam \lcount~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N11
dffeas \lcount[0] (
	.clk(!CLK),
	.d(\lcount~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(lcount[0]),
	.prn(vcc));
// synopsys translate_off
defparam \lcount[0] .is_wysiwyg = "true";
defparam \lcount[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N16
cycloneive_lcell_comb \lcount~3 (
// Equation(s):
// \lcount~3_combout  = (!\always0~3_combout  & (\Equal2~28_combout  & (lcount[0] $ (lcount[1]))))

	.dataa(lcount[0]),
	.datab(\always0~3_combout ),
	.datac(lcount[1]),
	.datad(\Equal2~28_combout ),
	.cin(gnd),
	.combout(\lcount~3_combout ),
	.cout());
// synopsys translate_off
defparam \lcount~3 .lut_mask = 16'h1200;
defparam \lcount~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N17
dffeas \lcount[1] (
	.clk(!CLK),
	.d(\lcount~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(lcount[1]),
	.prn(vcc));
// synopsys translate_off
defparam \lcount[1] .is_wysiwyg = "true";
defparam \lcount[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N22
cycloneive_lcell_comb \Add0~1 (
// Equation(s):
// \Add0~1_combout  = (lcount[2] $ (((!lcount[1]) # (!lcount[0])))) # (!\Equal2~28_combout )

	.dataa(lcount[0]),
	.datab(lcount[1]),
	.datac(lcount[2]),
	.datad(\Equal2~28_combout ),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~1 .lut_mask = 16'h87FF;
defparam \Add0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N8
cycloneive_lcell_comb \lcount~5 (
// Equation(s):
// \lcount~5_combout  = (!\always1~0_combout  & (!\always0~2_combout  & (!\Add0~1_combout  & \Equal2~28_combout )))

	.dataa(\always1~0_combout ),
	.datab(\always0~2_combout ),
	.datac(\Add0~1_combout ),
	.datad(\Equal2~28_combout ),
	.cin(gnd),
	.combout(\lcount~5_combout ),
	.cout());
// synopsys translate_off
defparam \lcount~5 .lut_mask = 16'h0100;
defparam \lcount~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N9
dffeas \lcount[2] (
	.clk(!CLK),
	.d(\lcount~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(lcount[2]),
	.prn(vcc));
// synopsys translate_off
defparam \lcount[2] .is_wysiwyg = "true";
defparam \lcount[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N20
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = (lcount[0] & (lcount[1] & (lcount[2] & \Equal2~28_combout )))

	.dataa(lcount[0]),
	.datab(lcount[1]),
	.datac(lcount[2]),
	.datad(\Equal2~28_combout ),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h8000;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N30
cycloneive_lcell_comb \lcount~2 (
// Equation(s):
// \lcount~2_combout  = (!\always0~3_combout  & (\Add0~0_combout  $ (((\Equal2~28_combout  & lcount[3])))))

	.dataa(\Equal2~28_combout ),
	.datab(\always0~3_combout ),
	.datac(lcount[3]),
	.datad(\Add0~0_combout ),
	.cin(gnd),
	.combout(\lcount~2_combout ),
	.cout());
// synopsys translate_off
defparam \lcount~2 .lut_mask = 16'h1320;
defparam \lcount~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N31
dffeas \lcount[3] (
	.clk(!CLK),
	.d(\lcount~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(lcount[3]),
	.prn(vcc));
// synopsys translate_off
defparam \lcount[3] .is_wysiwyg = "true";
defparam \lcount[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N28
cycloneive_lcell_comb \always1~1 (
// Equation(s):
// \always1~1_combout  = (lcount[3]) # ((lcount[2] & ((lcount[0]) # (lcount[1]))))

	.dataa(lcount[0]),
	.datab(lcount[3]),
	.datac(lcount[1]),
	.datad(lcount[2]),
	.cin(gnd),
	.combout(\always1~1_combout ),
	.cout());
// synopsys translate_off
defparam \always1~1 .lut_mask = 16'hFECC;
defparam \always1~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module altsyncram_1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramWEN,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramWEN;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



altsyncram_99f1 auto_generated(
	.ram_block3a32(ram_block3a32),
	.ram_block3a0(ram_block3a0),
	.ram_block3a33(ram_block3a33),
	.ram_block3a1(ram_block3a1),
	.ram_block3a34(ram_block3a34),
	.ram_block3a2(ram_block3a2),
	.ram_block3a35(ram_block3a35),
	.ram_block3a3(ram_block3a3),
	.ram_block3a36(ram_block3a36),
	.ram_block3a4(ram_block3a4),
	.ram_block3a37(ram_block3a37),
	.ram_block3a5(ram_block3a5),
	.ram_block3a38(ram_block3a38),
	.ram_block3a6(ram_block3a6),
	.ram_block3a39(ram_block3a39),
	.ram_block3a7(ram_block3a7),
	.ram_block3a40(ram_block3a40),
	.ram_block3a8(ram_block3a8),
	.ram_block3a41(ram_block3a41),
	.ram_block3a9(ram_block3a9),
	.ram_block3a42(ram_block3a42),
	.ram_block3a10(ram_block3a10),
	.ram_block3a43(ram_block3a43),
	.ram_block3a11(ram_block3a11),
	.ram_block3a44(ram_block3a44),
	.ram_block3a12(ram_block3a12),
	.ram_block3a45(ram_block3a45),
	.ram_block3a13(ram_block3a13),
	.ram_block3a46(ram_block3a46),
	.ram_block3a14(ram_block3a14),
	.ram_block3a47(ram_block3a47),
	.ram_block3a15(ram_block3a15),
	.ram_block3a48(ram_block3a48),
	.ram_block3a16(ram_block3a16),
	.ram_block3a49(ram_block3a49),
	.ram_block3a17(ram_block3a17),
	.ram_block3a50(ram_block3a50),
	.ram_block3a18(ram_block3a18),
	.ram_block3a51(ram_block3a51),
	.ram_block3a19(ram_block3a19),
	.ram_block3a52(ram_block3a52),
	.ram_block3a20(ram_block3a20),
	.ram_block3a53(ram_block3a53),
	.ram_block3a21(ram_block3a21),
	.ram_block3a54(ram_block3a54),
	.ram_block3a22(ram_block3a22),
	.ram_block3a55(ram_block3a55),
	.ram_block3a23(ram_block3a23),
	.ram_block3a56(ram_block3a56),
	.ram_block3a24(ram_block3a24),
	.ram_block3a57(ram_block3a57),
	.ram_block3a25(ram_block3a25),
	.ram_block3a58(ram_block3a58),
	.ram_block3a26(ram_block3a26),
	.ram_block3a59(ram_block3a59),
	.ram_block3a27(ram_block3a27),
	.ram_block3a60(ram_block3a60),
	.ram_block3a28(ram_block3a28),
	.ram_block3a61(ram_block3a61),
	.ram_block3a29(ram_block3a29),
	.ram_block3a62(ram_block3a62),
	.ram_block3a30(ram_block3a30),
	.ram_block3a63(ram_block3a63),
	.ram_block3a31(ram_block3a31),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.ramWEN(ramWEN),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.ramaddr1(ramaddr1),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_99f1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramWEN,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramWEN;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram1|ram_block3a32~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a0~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a33~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a1~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a34~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a2~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a35~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a3~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a36~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a4~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a37~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a5~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a38~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a6~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a39~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a7~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a40~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a8~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a41~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a9~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a42~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a10~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a43~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a11~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a44~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a12~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a45~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a13~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a46~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a14~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a47~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a15~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a48~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a16~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a49~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a17~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a50~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a18~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a51~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a19~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a52~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a20~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a53~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a21~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a54~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a22~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a55~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a23~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a56~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a24~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a57~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a25~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a58~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a26~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a59~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a27~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a60~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a28~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a61~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a29~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a62~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a30~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a63~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a31~PORTBDATAOUT0 ;
wire \mgl_prim2|sdr~0_combout ;
wire [0:0] \altsyncram1|address_reg_b ;
wire [31:0] \mgl_prim2|ram_rom_data_reg ;
wire [13:0] \mgl_prim2|ram_rom_addr_reg ;


sld_mod_ram_rom mgl_prim2(
	.ram_block3a32(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a0(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a33(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a1(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a34(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a2(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a35(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a3(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a36(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a4(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a37(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a5(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a38(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a6(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a39(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a7(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a40(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a8(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a41(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a9(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a42(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a10(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a43(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a11(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a44(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a12(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a45(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a13(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a46(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a14(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a47(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a15(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a48(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a16(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a49(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a17(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a50(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a18(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a51(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a19(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a52(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a20(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a53(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a21(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a54(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a22(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a55(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a23(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a56(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a24(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a57(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a25(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a58(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a26(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a59(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a27(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a60(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a28(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a61(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a29(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a62(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a30(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a63(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a31(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.is_in_use_reg1(is_in_use_reg),
	.ram_rom_data_reg_0(\mgl_prim2|ram_rom_data_reg [0]),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.ram_rom_addr_reg_0(\mgl_prim2|ram_rom_addr_reg [0]),
	.ram_rom_addr_reg_1(\mgl_prim2|ram_rom_addr_reg [1]),
	.ram_rom_addr_reg_2(\mgl_prim2|ram_rom_addr_reg [2]),
	.ram_rom_addr_reg_3(\mgl_prim2|ram_rom_addr_reg [3]),
	.ram_rom_addr_reg_4(\mgl_prim2|ram_rom_addr_reg [4]),
	.ram_rom_addr_reg_5(\mgl_prim2|ram_rom_addr_reg [5]),
	.ram_rom_addr_reg_6(\mgl_prim2|ram_rom_addr_reg [6]),
	.ram_rom_addr_reg_7(\mgl_prim2|ram_rom_addr_reg [7]),
	.ram_rom_addr_reg_8(\mgl_prim2|ram_rom_addr_reg [8]),
	.ram_rom_addr_reg_9(\mgl_prim2|ram_rom_addr_reg [9]),
	.ram_rom_addr_reg_10(\mgl_prim2|ram_rom_addr_reg [10]),
	.ram_rom_addr_reg_11(\mgl_prim2|ram_rom_addr_reg [11]),
	.ram_rom_addr_reg_12(\mgl_prim2|ram_rom_addr_reg [12]),
	.ram_rom_data_reg_1(\mgl_prim2|ram_rom_data_reg [1]),
	.ram_rom_data_reg_2(\mgl_prim2|ram_rom_data_reg [2]),
	.ram_rom_data_reg_3(\mgl_prim2|ram_rom_data_reg [3]),
	.ram_rom_data_reg_4(\mgl_prim2|ram_rom_data_reg [4]),
	.ram_rom_data_reg_5(\mgl_prim2|ram_rom_data_reg [5]),
	.ram_rom_data_reg_6(\mgl_prim2|ram_rom_data_reg [6]),
	.ram_rom_data_reg_7(\mgl_prim2|ram_rom_data_reg [7]),
	.ram_rom_data_reg_8(\mgl_prim2|ram_rom_data_reg [8]),
	.ram_rom_data_reg_9(\mgl_prim2|ram_rom_data_reg [9]),
	.ram_rom_data_reg_10(\mgl_prim2|ram_rom_data_reg [10]),
	.ram_rom_data_reg_11(\mgl_prim2|ram_rom_data_reg [11]),
	.ram_rom_data_reg_12(\mgl_prim2|ram_rom_data_reg [12]),
	.ram_rom_data_reg_13(\mgl_prim2|ram_rom_data_reg [13]),
	.ram_rom_data_reg_14(\mgl_prim2|ram_rom_data_reg [14]),
	.ram_rom_data_reg_15(\mgl_prim2|ram_rom_data_reg [15]),
	.ram_rom_data_reg_16(\mgl_prim2|ram_rom_data_reg [16]),
	.ram_rom_data_reg_17(\mgl_prim2|ram_rom_data_reg [17]),
	.ram_rom_data_reg_18(\mgl_prim2|ram_rom_data_reg [18]),
	.ram_rom_data_reg_19(\mgl_prim2|ram_rom_data_reg [19]),
	.ram_rom_data_reg_20(\mgl_prim2|ram_rom_data_reg [20]),
	.ram_rom_data_reg_21(\mgl_prim2|ram_rom_data_reg [21]),
	.ram_rom_data_reg_22(\mgl_prim2|ram_rom_data_reg [22]),
	.ram_rom_data_reg_23(\mgl_prim2|ram_rom_data_reg [23]),
	.ram_rom_data_reg_24(\mgl_prim2|ram_rom_data_reg [24]),
	.ram_rom_data_reg_25(\mgl_prim2|ram_rom_data_reg [25]),
	.ram_rom_data_reg_26(\mgl_prim2|ram_rom_data_reg [26]),
	.ram_rom_data_reg_27(\mgl_prim2|ram_rom_data_reg [27]),
	.ram_rom_data_reg_28(\mgl_prim2|ram_rom_data_reg [28]),
	.ram_rom_data_reg_29(\mgl_prim2|ram_rom_data_reg [29]),
	.ram_rom_data_reg_30(\mgl_prim2|ram_rom_data_reg [30]),
	.ram_rom_data_reg_31(\mgl_prim2|ram_rom_data_reg [31]),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.ir_in({gnd,irf_reg_3_1,gnd,gnd,irf_reg_0_1}),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.raw_tck(altera_internal_jtag1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

altsyncram_fta2 altsyncram1(
	.ram_block3a321(ram_block3a32),
	.ram_block3a322(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a01(ram_block3a0),
	.ram_block3a02(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a331(ram_block3a33),
	.ram_block3a332(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a110(ram_block3a1),
	.ram_block3a111(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a341(ram_block3a34),
	.ram_block3a342(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a210(ram_block3a2),
	.ram_block3a211(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a351(ram_block3a35),
	.ram_block3a352(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a310(ram_block3a3),
	.ram_block3a311(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a361(ram_block3a36),
	.ram_block3a362(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a410(ram_block3a4),
	.ram_block3a411(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a371(ram_block3a37),
	.ram_block3a372(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a510(ram_block3a5),
	.ram_block3a511(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a381(ram_block3a38),
	.ram_block3a382(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a64(ram_block3a6),
	.ram_block3a65(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a391(ram_block3a39),
	.ram_block3a392(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a71(ram_block3a7),
	.ram_block3a72(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a401(ram_block3a40),
	.ram_block3a402(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a81(ram_block3a8),
	.ram_block3a82(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a412(ram_block3a41),
	.ram_block3a413(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a91(ram_block3a9),
	.ram_block3a92(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a421(ram_block3a42),
	.ram_block3a422(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a101(ram_block3a10),
	.ram_block3a102(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a431(ram_block3a43),
	.ram_block3a432(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a112(ram_block3a11),
	.ram_block3a113(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a441(ram_block3a44),
	.ram_block3a442(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a121(ram_block3a12),
	.ram_block3a122(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a451(ram_block3a45),
	.ram_block3a452(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a131(ram_block3a13),
	.ram_block3a132(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a461(ram_block3a46),
	.ram_block3a462(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a141(ram_block3a14),
	.ram_block3a142(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a471(ram_block3a47),
	.ram_block3a472(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a151(ram_block3a15),
	.ram_block3a152(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a481(ram_block3a48),
	.ram_block3a482(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a161(ram_block3a16),
	.ram_block3a162(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a491(ram_block3a49),
	.ram_block3a492(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a171(ram_block3a17),
	.ram_block3a172(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a501(ram_block3a50),
	.ram_block3a502(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a181(ram_block3a18),
	.ram_block3a182(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a512(ram_block3a51),
	.ram_block3a513(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a191(ram_block3a19),
	.ram_block3a192(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a521(ram_block3a52),
	.ram_block3a522(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a201(ram_block3a20),
	.ram_block3a202(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a531(ram_block3a53),
	.ram_block3a532(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a212(ram_block3a21),
	.ram_block3a213(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a541(ram_block3a54),
	.ram_block3a542(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a221(ram_block3a22),
	.ram_block3a222(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a551(ram_block3a55),
	.ram_block3a552(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a231(ram_block3a23),
	.ram_block3a232(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a561(ram_block3a56),
	.ram_block3a562(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a241(ram_block3a24),
	.ram_block3a242(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a571(ram_block3a57),
	.ram_block3a572(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a251(ram_block3a25),
	.ram_block3a252(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a581(ram_block3a58),
	.ram_block3a582(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a261(ram_block3a26),
	.ram_block3a262(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a591(ram_block3a59),
	.ram_block3a592(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a271(ram_block3a27),
	.ram_block3a272(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a601(ram_block3a60),
	.ram_block3a602(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a281(ram_block3a28),
	.ram_block3a282(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a611(ram_block3a61),
	.ram_block3a612(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a291(ram_block3a29),
	.ram_block3a292(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a621(ram_block3a62),
	.ram_block3a622(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a301(ram_block3a30),
	.ram_block3a302(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a631(ram_block3a63),
	.ram_block3a632(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a312(ram_block3a31),
	.ram_block3a313(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.data_b({\mgl_prim2|ram_rom_data_reg [31],\mgl_prim2|ram_rom_data_reg [30],\mgl_prim2|ram_rom_data_reg [29],\mgl_prim2|ram_rom_data_reg [28],\mgl_prim2|ram_rom_data_reg [27],\mgl_prim2|ram_rom_data_reg [26],\mgl_prim2|ram_rom_data_reg [25],\mgl_prim2|ram_rom_data_reg [24],\mgl_prim2|ram_rom_data_reg [23],
\mgl_prim2|ram_rom_data_reg [22],\mgl_prim2|ram_rom_data_reg [21],\mgl_prim2|ram_rom_data_reg [20],\mgl_prim2|ram_rom_data_reg [19],\mgl_prim2|ram_rom_data_reg [18],\mgl_prim2|ram_rom_data_reg [17],\mgl_prim2|ram_rom_data_reg [16],\mgl_prim2|ram_rom_data_reg [15],\mgl_prim2|ram_rom_data_reg [14],
\mgl_prim2|ram_rom_data_reg [13],\mgl_prim2|ram_rom_data_reg [12],\mgl_prim2|ram_rom_data_reg [11],\mgl_prim2|ram_rom_data_reg [10],\mgl_prim2|ram_rom_data_reg [9],\mgl_prim2|ram_rom_data_reg [8],\mgl_prim2|ram_rom_data_reg [7],\mgl_prim2|ram_rom_data_reg [6],\mgl_prim2|ram_rom_data_reg [5],
\mgl_prim2|ram_rom_data_reg [4],\mgl_prim2|ram_rom_data_reg [3],\mgl_prim2|ram_rom_data_reg [2],\mgl_prim2|ram_rom_data_reg [1],\mgl_prim2|ram_rom_data_reg [0]}),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.address_b({gnd,\mgl_prim2|ram_rom_addr_reg [12],\mgl_prim2|ram_rom_addr_reg [11],\mgl_prim2|ram_rom_addr_reg [10],\mgl_prim2|ram_rom_addr_reg [9],\mgl_prim2|ram_rom_addr_reg [8],\mgl_prim2|ram_rom_addr_reg [7],\mgl_prim2|ram_rom_addr_reg [6],\mgl_prim2|ram_rom_addr_reg [5],\mgl_prim2|ram_rom_addr_reg [4],
\mgl_prim2|ram_rom_addr_reg [3],\mgl_prim2|ram_rom_addr_reg [2],\mgl_prim2|ram_rom_addr_reg [1],\mgl_prim2|ram_rom_addr_reg [0]}),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.always1(always1),
	.ramWEN(ramWEN),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.ramaddr1(ramaddr1),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.clock1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_fta2 (
	ram_block3a321,
	ram_block3a322,
	ram_block3a01,
	ram_block3a02,
	ram_block3a331,
	ram_block3a332,
	ram_block3a110,
	ram_block3a111,
	ram_block3a341,
	ram_block3a342,
	ram_block3a210,
	ram_block3a211,
	ram_block3a351,
	ram_block3a352,
	ram_block3a310,
	ram_block3a311,
	ram_block3a361,
	ram_block3a362,
	ram_block3a410,
	ram_block3a411,
	ram_block3a371,
	ram_block3a372,
	ram_block3a510,
	ram_block3a511,
	ram_block3a381,
	ram_block3a382,
	ram_block3a64,
	ram_block3a65,
	ram_block3a391,
	ram_block3a392,
	ram_block3a71,
	ram_block3a72,
	ram_block3a401,
	ram_block3a402,
	ram_block3a81,
	ram_block3a82,
	ram_block3a412,
	ram_block3a413,
	ram_block3a91,
	ram_block3a92,
	ram_block3a421,
	ram_block3a422,
	ram_block3a101,
	ram_block3a102,
	ram_block3a431,
	ram_block3a432,
	ram_block3a112,
	ram_block3a113,
	ram_block3a441,
	ram_block3a442,
	ram_block3a121,
	ram_block3a122,
	ram_block3a451,
	ram_block3a452,
	ram_block3a131,
	ram_block3a132,
	ram_block3a461,
	ram_block3a462,
	ram_block3a141,
	ram_block3a142,
	ram_block3a471,
	ram_block3a472,
	ram_block3a151,
	ram_block3a152,
	ram_block3a481,
	ram_block3a482,
	ram_block3a161,
	ram_block3a162,
	ram_block3a491,
	ram_block3a492,
	ram_block3a171,
	ram_block3a172,
	ram_block3a501,
	ram_block3a502,
	ram_block3a181,
	ram_block3a182,
	ram_block3a512,
	ram_block3a513,
	ram_block3a191,
	ram_block3a192,
	ram_block3a521,
	ram_block3a522,
	ram_block3a201,
	ram_block3a202,
	ram_block3a531,
	ram_block3a532,
	ram_block3a212,
	ram_block3a213,
	ram_block3a541,
	ram_block3a542,
	ram_block3a221,
	ram_block3a222,
	ram_block3a551,
	ram_block3a552,
	ram_block3a231,
	ram_block3a232,
	ram_block3a561,
	ram_block3a562,
	ram_block3a241,
	ram_block3a242,
	ram_block3a571,
	ram_block3a572,
	ram_block3a251,
	ram_block3a252,
	ram_block3a581,
	ram_block3a582,
	ram_block3a261,
	ram_block3a262,
	ram_block3a591,
	ram_block3a592,
	ram_block3a271,
	ram_block3a272,
	ram_block3a601,
	ram_block3a602,
	ram_block3a281,
	ram_block3a282,
	ram_block3a611,
	ram_block3a612,
	ram_block3a291,
	ram_block3a292,
	ram_block3a621,
	ram_block3a622,
	ram_block3a301,
	ram_block3a302,
	ram_block3a631,
	ram_block3a632,
	ram_block3a312,
	ram_block3a313,
	data_b,
	ram_rom_addr_reg_13,
	address_b,
	address_reg_a_0,
	address_a,
	ramaddr,
	always1,
	ramWEN,
	sdr,
	data_a,
	address_reg_b_0,
	ramaddr1,
	irf_reg_2_1,
	state_5,
	clock1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a321;
output 	ram_block3a322;
output 	ram_block3a01;
output 	ram_block3a02;
output 	ram_block3a331;
output 	ram_block3a332;
output 	ram_block3a110;
output 	ram_block3a111;
output 	ram_block3a341;
output 	ram_block3a342;
output 	ram_block3a210;
output 	ram_block3a211;
output 	ram_block3a351;
output 	ram_block3a352;
output 	ram_block3a310;
output 	ram_block3a311;
output 	ram_block3a361;
output 	ram_block3a362;
output 	ram_block3a410;
output 	ram_block3a411;
output 	ram_block3a371;
output 	ram_block3a372;
output 	ram_block3a510;
output 	ram_block3a511;
output 	ram_block3a381;
output 	ram_block3a382;
output 	ram_block3a64;
output 	ram_block3a65;
output 	ram_block3a391;
output 	ram_block3a392;
output 	ram_block3a71;
output 	ram_block3a72;
output 	ram_block3a401;
output 	ram_block3a402;
output 	ram_block3a81;
output 	ram_block3a82;
output 	ram_block3a412;
output 	ram_block3a413;
output 	ram_block3a91;
output 	ram_block3a92;
output 	ram_block3a421;
output 	ram_block3a422;
output 	ram_block3a101;
output 	ram_block3a102;
output 	ram_block3a431;
output 	ram_block3a432;
output 	ram_block3a112;
output 	ram_block3a113;
output 	ram_block3a441;
output 	ram_block3a442;
output 	ram_block3a121;
output 	ram_block3a122;
output 	ram_block3a451;
output 	ram_block3a452;
output 	ram_block3a131;
output 	ram_block3a132;
output 	ram_block3a461;
output 	ram_block3a462;
output 	ram_block3a141;
output 	ram_block3a142;
output 	ram_block3a471;
output 	ram_block3a472;
output 	ram_block3a151;
output 	ram_block3a152;
output 	ram_block3a481;
output 	ram_block3a482;
output 	ram_block3a161;
output 	ram_block3a162;
output 	ram_block3a491;
output 	ram_block3a492;
output 	ram_block3a171;
output 	ram_block3a172;
output 	ram_block3a501;
output 	ram_block3a502;
output 	ram_block3a181;
output 	ram_block3a182;
output 	ram_block3a512;
output 	ram_block3a513;
output 	ram_block3a191;
output 	ram_block3a192;
output 	ram_block3a521;
output 	ram_block3a522;
output 	ram_block3a201;
output 	ram_block3a202;
output 	ram_block3a531;
output 	ram_block3a532;
output 	ram_block3a212;
output 	ram_block3a213;
output 	ram_block3a541;
output 	ram_block3a542;
output 	ram_block3a221;
output 	ram_block3a222;
output 	ram_block3a551;
output 	ram_block3a552;
output 	ram_block3a231;
output 	ram_block3a232;
output 	ram_block3a561;
output 	ram_block3a562;
output 	ram_block3a241;
output 	ram_block3a242;
output 	ram_block3a571;
output 	ram_block3a572;
output 	ram_block3a251;
output 	ram_block3a252;
output 	ram_block3a581;
output 	ram_block3a582;
output 	ram_block3a261;
output 	ram_block3a262;
output 	ram_block3a591;
output 	ram_block3a592;
output 	ram_block3a271;
output 	ram_block3a272;
output 	ram_block3a601;
output 	ram_block3a602;
output 	ram_block3a281;
output 	ram_block3a282;
output 	ram_block3a611;
output 	ram_block3a612;
output 	ram_block3a291;
output 	ram_block3a292;
output 	ram_block3a621;
output 	ram_block3a622;
output 	ram_block3a301;
output 	ram_block3a302;
output 	ram_block3a631;
output 	ram_block3a632;
output 	ram_block3a312;
output 	ram_block3a313;
input 	[31:0] data_b;
input 	ram_rom_addr_reg_13;
input 	[13:0] address_b;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	always1;
input 	ramWEN;
input 	sdr;
input 	[31:0] data_a;
output 	address_reg_b_0;
input 	ramaddr1;
input 	irf_reg_2_1;
input 	state_5;
input 	clock1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \decode4|eq_node[1]~0_combout ;
wire \decode5|eq_node[1]~0_combout ;
wire \decode4|eq_node[0]~1_combout ;
wire \decode5|eq_node[0]~1_combout ;
wire \address_reg_b[0]~feeder_combout ;

wire [0:0] ram_block3a32_PORTADATAOUT_bus;
wire [0:0] ram_block3a32_PORTBDATAOUT_bus;
wire [0:0] ram_block3a0_PORTADATAOUT_bus;
wire [0:0] ram_block3a0_PORTBDATAOUT_bus;
wire [0:0] ram_block3a33_PORTADATAOUT_bus;
wire [0:0] ram_block3a33_PORTBDATAOUT_bus;
wire [0:0] ram_block3a1_PORTADATAOUT_bus;
wire [0:0] ram_block3a1_PORTBDATAOUT_bus;
wire [0:0] ram_block3a34_PORTADATAOUT_bus;
wire [0:0] ram_block3a34_PORTBDATAOUT_bus;
wire [0:0] ram_block3a2_PORTADATAOUT_bus;
wire [0:0] ram_block3a2_PORTBDATAOUT_bus;
wire [0:0] ram_block3a35_PORTADATAOUT_bus;
wire [0:0] ram_block3a35_PORTBDATAOUT_bus;
wire [0:0] ram_block3a3_PORTADATAOUT_bus;
wire [0:0] ram_block3a3_PORTBDATAOUT_bus;
wire [0:0] ram_block3a36_PORTADATAOUT_bus;
wire [0:0] ram_block3a36_PORTBDATAOUT_bus;
wire [0:0] ram_block3a4_PORTADATAOUT_bus;
wire [0:0] ram_block3a4_PORTBDATAOUT_bus;
wire [0:0] ram_block3a37_PORTADATAOUT_bus;
wire [0:0] ram_block3a37_PORTBDATAOUT_bus;
wire [0:0] ram_block3a5_PORTADATAOUT_bus;
wire [0:0] ram_block3a5_PORTBDATAOUT_bus;
wire [0:0] ram_block3a38_PORTADATAOUT_bus;
wire [0:0] ram_block3a38_PORTBDATAOUT_bus;
wire [0:0] ram_block3a6_PORTADATAOUT_bus;
wire [0:0] ram_block3a6_PORTBDATAOUT_bus;
wire [0:0] ram_block3a39_PORTADATAOUT_bus;
wire [0:0] ram_block3a39_PORTBDATAOUT_bus;
wire [0:0] ram_block3a7_PORTADATAOUT_bus;
wire [0:0] ram_block3a7_PORTBDATAOUT_bus;
wire [0:0] ram_block3a40_PORTADATAOUT_bus;
wire [0:0] ram_block3a40_PORTBDATAOUT_bus;
wire [0:0] ram_block3a8_PORTADATAOUT_bus;
wire [0:0] ram_block3a8_PORTBDATAOUT_bus;
wire [0:0] ram_block3a41_PORTADATAOUT_bus;
wire [0:0] ram_block3a41_PORTBDATAOUT_bus;
wire [0:0] ram_block3a9_PORTADATAOUT_bus;
wire [0:0] ram_block3a9_PORTBDATAOUT_bus;
wire [0:0] ram_block3a42_PORTADATAOUT_bus;
wire [0:0] ram_block3a42_PORTBDATAOUT_bus;
wire [0:0] ram_block3a10_PORTADATAOUT_bus;
wire [0:0] ram_block3a10_PORTBDATAOUT_bus;
wire [0:0] ram_block3a43_PORTADATAOUT_bus;
wire [0:0] ram_block3a43_PORTBDATAOUT_bus;
wire [0:0] ram_block3a11_PORTADATAOUT_bus;
wire [0:0] ram_block3a11_PORTBDATAOUT_bus;
wire [0:0] ram_block3a44_PORTADATAOUT_bus;
wire [0:0] ram_block3a44_PORTBDATAOUT_bus;
wire [0:0] ram_block3a12_PORTADATAOUT_bus;
wire [0:0] ram_block3a12_PORTBDATAOUT_bus;
wire [0:0] ram_block3a45_PORTADATAOUT_bus;
wire [0:0] ram_block3a45_PORTBDATAOUT_bus;
wire [0:0] ram_block3a13_PORTADATAOUT_bus;
wire [0:0] ram_block3a13_PORTBDATAOUT_bus;
wire [0:0] ram_block3a46_PORTADATAOUT_bus;
wire [0:0] ram_block3a46_PORTBDATAOUT_bus;
wire [0:0] ram_block3a14_PORTADATAOUT_bus;
wire [0:0] ram_block3a14_PORTBDATAOUT_bus;
wire [0:0] ram_block3a47_PORTADATAOUT_bus;
wire [0:0] ram_block3a47_PORTBDATAOUT_bus;
wire [0:0] ram_block3a15_PORTADATAOUT_bus;
wire [0:0] ram_block3a15_PORTBDATAOUT_bus;
wire [0:0] ram_block3a48_PORTADATAOUT_bus;
wire [0:0] ram_block3a48_PORTBDATAOUT_bus;
wire [0:0] ram_block3a16_PORTADATAOUT_bus;
wire [0:0] ram_block3a16_PORTBDATAOUT_bus;
wire [0:0] ram_block3a49_PORTADATAOUT_bus;
wire [0:0] ram_block3a49_PORTBDATAOUT_bus;
wire [0:0] ram_block3a17_PORTADATAOUT_bus;
wire [0:0] ram_block3a17_PORTBDATAOUT_bus;
wire [0:0] ram_block3a50_PORTADATAOUT_bus;
wire [0:0] ram_block3a50_PORTBDATAOUT_bus;
wire [0:0] ram_block3a18_PORTADATAOUT_bus;
wire [0:0] ram_block3a18_PORTBDATAOUT_bus;
wire [0:0] ram_block3a51_PORTADATAOUT_bus;
wire [0:0] ram_block3a51_PORTBDATAOUT_bus;
wire [0:0] ram_block3a19_PORTADATAOUT_bus;
wire [0:0] ram_block3a19_PORTBDATAOUT_bus;
wire [0:0] ram_block3a52_PORTADATAOUT_bus;
wire [0:0] ram_block3a52_PORTBDATAOUT_bus;
wire [0:0] ram_block3a20_PORTADATAOUT_bus;
wire [0:0] ram_block3a20_PORTBDATAOUT_bus;
wire [0:0] ram_block3a53_PORTADATAOUT_bus;
wire [0:0] ram_block3a53_PORTBDATAOUT_bus;
wire [0:0] ram_block3a21_PORTADATAOUT_bus;
wire [0:0] ram_block3a21_PORTBDATAOUT_bus;
wire [0:0] ram_block3a54_PORTADATAOUT_bus;
wire [0:0] ram_block3a54_PORTBDATAOUT_bus;
wire [0:0] ram_block3a22_PORTADATAOUT_bus;
wire [0:0] ram_block3a22_PORTBDATAOUT_bus;
wire [0:0] ram_block3a55_PORTADATAOUT_bus;
wire [0:0] ram_block3a55_PORTBDATAOUT_bus;
wire [0:0] ram_block3a23_PORTADATAOUT_bus;
wire [0:0] ram_block3a23_PORTBDATAOUT_bus;
wire [0:0] ram_block3a56_PORTADATAOUT_bus;
wire [0:0] ram_block3a56_PORTBDATAOUT_bus;
wire [0:0] ram_block3a24_PORTADATAOUT_bus;
wire [0:0] ram_block3a24_PORTBDATAOUT_bus;
wire [0:0] ram_block3a57_PORTADATAOUT_bus;
wire [0:0] ram_block3a57_PORTBDATAOUT_bus;
wire [0:0] ram_block3a25_PORTADATAOUT_bus;
wire [0:0] ram_block3a25_PORTBDATAOUT_bus;
wire [0:0] ram_block3a58_PORTADATAOUT_bus;
wire [0:0] ram_block3a58_PORTBDATAOUT_bus;
wire [0:0] ram_block3a26_PORTADATAOUT_bus;
wire [0:0] ram_block3a26_PORTBDATAOUT_bus;
wire [0:0] ram_block3a59_PORTADATAOUT_bus;
wire [0:0] ram_block3a59_PORTBDATAOUT_bus;
wire [0:0] ram_block3a27_PORTADATAOUT_bus;
wire [0:0] ram_block3a27_PORTBDATAOUT_bus;
wire [0:0] ram_block3a60_PORTADATAOUT_bus;
wire [0:0] ram_block3a60_PORTBDATAOUT_bus;
wire [0:0] ram_block3a28_PORTADATAOUT_bus;
wire [0:0] ram_block3a28_PORTBDATAOUT_bus;
wire [0:0] ram_block3a61_PORTADATAOUT_bus;
wire [0:0] ram_block3a61_PORTBDATAOUT_bus;
wire [0:0] ram_block3a29_PORTADATAOUT_bus;
wire [0:0] ram_block3a29_PORTBDATAOUT_bus;
wire [0:0] ram_block3a62_PORTADATAOUT_bus;
wire [0:0] ram_block3a62_PORTBDATAOUT_bus;
wire [0:0] ram_block3a30_PORTADATAOUT_bus;
wire [0:0] ram_block3a30_PORTBDATAOUT_bus;
wire [0:0] ram_block3a63_PORTADATAOUT_bus;
wire [0:0] ram_block3a63_PORTBDATAOUT_bus;
wire [0:0] ram_block3a31_PORTADATAOUT_bus;
wire [0:0] ram_block3a31_PORTBDATAOUT_bus;

assign ram_block3a321 = ram_block3a32_PORTADATAOUT_bus[0];

assign ram_block3a322 = ram_block3a32_PORTBDATAOUT_bus[0];

assign ram_block3a01 = ram_block3a0_PORTADATAOUT_bus[0];

assign ram_block3a02 = ram_block3a0_PORTBDATAOUT_bus[0];

assign ram_block3a331 = ram_block3a33_PORTADATAOUT_bus[0];

assign ram_block3a332 = ram_block3a33_PORTBDATAOUT_bus[0];

assign ram_block3a110 = ram_block3a1_PORTADATAOUT_bus[0];

assign ram_block3a111 = ram_block3a1_PORTBDATAOUT_bus[0];

assign ram_block3a341 = ram_block3a34_PORTADATAOUT_bus[0];

assign ram_block3a342 = ram_block3a34_PORTBDATAOUT_bus[0];

assign ram_block3a210 = ram_block3a2_PORTADATAOUT_bus[0];

assign ram_block3a211 = ram_block3a2_PORTBDATAOUT_bus[0];

assign ram_block3a351 = ram_block3a35_PORTADATAOUT_bus[0];

assign ram_block3a352 = ram_block3a35_PORTBDATAOUT_bus[0];

assign ram_block3a310 = ram_block3a3_PORTADATAOUT_bus[0];

assign ram_block3a311 = ram_block3a3_PORTBDATAOUT_bus[0];

assign ram_block3a361 = ram_block3a36_PORTADATAOUT_bus[0];

assign ram_block3a362 = ram_block3a36_PORTBDATAOUT_bus[0];

assign ram_block3a410 = ram_block3a4_PORTADATAOUT_bus[0];

assign ram_block3a411 = ram_block3a4_PORTBDATAOUT_bus[0];

assign ram_block3a371 = ram_block3a37_PORTADATAOUT_bus[0];

assign ram_block3a372 = ram_block3a37_PORTBDATAOUT_bus[0];

assign ram_block3a510 = ram_block3a5_PORTADATAOUT_bus[0];

assign ram_block3a511 = ram_block3a5_PORTBDATAOUT_bus[0];

assign ram_block3a381 = ram_block3a38_PORTADATAOUT_bus[0];

assign ram_block3a382 = ram_block3a38_PORTBDATAOUT_bus[0];

assign ram_block3a64 = ram_block3a6_PORTADATAOUT_bus[0];

assign ram_block3a65 = ram_block3a6_PORTBDATAOUT_bus[0];

assign ram_block3a391 = ram_block3a39_PORTADATAOUT_bus[0];

assign ram_block3a392 = ram_block3a39_PORTBDATAOUT_bus[0];

assign ram_block3a71 = ram_block3a7_PORTADATAOUT_bus[0];

assign ram_block3a72 = ram_block3a7_PORTBDATAOUT_bus[0];

assign ram_block3a401 = ram_block3a40_PORTADATAOUT_bus[0];

assign ram_block3a402 = ram_block3a40_PORTBDATAOUT_bus[0];

assign ram_block3a81 = ram_block3a8_PORTADATAOUT_bus[0];

assign ram_block3a82 = ram_block3a8_PORTBDATAOUT_bus[0];

assign ram_block3a412 = ram_block3a41_PORTADATAOUT_bus[0];

assign ram_block3a413 = ram_block3a41_PORTBDATAOUT_bus[0];

assign ram_block3a91 = ram_block3a9_PORTADATAOUT_bus[0];

assign ram_block3a92 = ram_block3a9_PORTBDATAOUT_bus[0];

assign ram_block3a421 = ram_block3a42_PORTADATAOUT_bus[0];

assign ram_block3a422 = ram_block3a42_PORTBDATAOUT_bus[0];

assign ram_block3a101 = ram_block3a10_PORTADATAOUT_bus[0];

assign ram_block3a102 = ram_block3a10_PORTBDATAOUT_bus[0];

assign ram_block3a431 = ram_block3a43_PORTADATAOUT_bus[0];

assign ram_block3a432 = ram_block3a43_PORTBDATAOUT_bus[0];

assign ram_block3a112 = ram_block3a11_PORTADATAOUT_bus[0];

assign ram_block3a113 = ram_block3a11_PORTBDATAOUT_bus[0];

assign ram_block3a441 = ram_block3a44_PORTADATAOUT_bus[0];

assign ram_block3a442 = ram_block3a44_PORTBDATAOUT_bus[0];

assign ram_block3a121 = ram_block3a12_PORTADATAOUT_bus[0];

assign ram_block3a122 = ram_block3a12_PORTBDATAOUT_bus[0];

assign ram_block3a451 = ram_block3a45_PORTADATAOUT_bus[0];

assign ram_block3a452 = ram_block3a45_PORTBDATAOUT_bus[0];

assign ram_block3a131 = ram_block3a13_PORTADATAOUT_bus[0];

assign ram_block3a132 = ram_block3a13_PORTBDATAOUT_bus[0];

assign ram_block3a461 = ram_block3a46_PORTADATAOUT_bus[0];

assign ram_block3a462 = ram_block3a46_PORTBDATAOUT_bus[0];

assign ram_block3a141 = ram_block3a14_PORTADATAOUT_bus[0];

assign ram_block3a142 = ram_block3a14_PORTBDATAOUT_bus[0];

assign ram_block3a471 = ram_block3a47_PORTADATAOUT_bus[0];

assign ram_block3a472 = ram_block3a47_PORTBDATAOUT_bus[0];

assign ram_block3a151 = ram_block3a15_PORTADATAOUT_bus[0];

assign ram_block3a152 = ram_block3a15_PORTBDATAOUT_bus[0];

assign ram_block3a481 = ram_block3a48_PORTADATAOUT_bus[0];

assign ram_block3a482 = ram_block3a48_PORTBDATAOUT_bus[0];

assign ram_block3a161 = ram_block3a16_PORTADATAOUT_bus[0];

assign ram_block3a162 = ram_block3a16_PORTBDATAOUT_bus[0];

assign ram_block3a491 = ram_block3a49_PORTADATAOUT_bus[0];

assign ram_block3a492 = ram_block3a49_PORTBDATAOUT_bus[0];

assign ram_block3a171 = ram_block3a17_PORTADATAOUT_bus[0];

assign ram_block3a172 = ram_block3a17_PORTBDATAOUT_bus[0];

assign ram_block3a501 = ram_block3a50_PORTADATAOUT_bus[0];

assign ram_block3a502 = ram_block3a50_PORTBDATAOUT_bus[0];

assign ram_block3a181 = ram_block3a18_PORTADATAOUT_bus[0];

assign ram_block3a182 = ram_block3a18_PORTBDATAOUT_bus[0];

assign ram_block3a512 = ram_block3a51_PORTADATAOUT_bus[0];

assign ram_block3a513 = ram_block3a51_PORTBDATAOUT_bus[0];

assign ram_block3a191 = ram_block3a19_PORTADATAOUT_bus[0];

assign ram_block3a192 = ram_block3a19_PORTBDATAOUT_bus[0];

assign ram_block3a521 = ram_block3a52_PORTADATAOUT_bus[0];

assign ram_block3a522 = ram_block3a52_PORTBDATAOUT_bus[0];

assign ram_block3a201 = ram_block3a20_PORTADATAOUT_bus[0];

assign ram_block3a202 = ram_block3a20_PORTBDATAOUT_bus[0];

assign ram_block3a531 = ram_block3a53_PORTADATAOUT_bus[0];

assign ram_block3a532 = ram_block3a53_PORTBDATAOUT_bus[0];

assign ram_block3a212 = ram_block3a21_PORTADATAOUT_bus[0];

assign ram_block3a213 = ram_block3a21_PORTBDATAOUT_bus[0];

assign ram_block3a541 = ram_block3a54_PORTADATAOUT_bus[0];

assign ram_block3a542 = ram_block3a54_PORTBDATAOUT_bus[0];

assign ram_block3a221 = ram_block3a22_PORTADATAOUT_bus[0];

assign ram_block3a222 = ram_block3a22_PORTBDATAOUT_bus[0];

assign ram_block3a551 = ram_block3a55_PORTADATAOUT_bus[0];

assign ram_block3a552 = ram_block3a55_PORTBDATAOUT_bus[0];

assign ram_block3a231 = ram_block3a23_PORTADATAOUT_bus[0];

assign ram_block3a232 = ram_block3a23_PORTBDATAOUT_bus[0];

assign ram_block3a561 = ram_block3a56_PORTADATAOUT_bus[0];

assign ram_block3a562 = ram_block3a56_PORTBDATAOUT_bus[0];

assign ram_block3a241 = ram_block3a24_PORTADATAOUT_bus[0];

assign ram_block3a242 = ram_block3a24_PORTBDATAOUT_bus[0];

assign ram_block3a571 = ram_block3a57_PORTADATAOUT_bus[0];

assign ram_block3a572 = ram_block3a57_PORTBDATAOUT_bus[0];

assign ram_block3a251 = ram_block3a25_PORTADATAOUT_bus[0];

assign ram_block3a252 = ram_block3a25_PORTBDATAOUT_bus[0];

assign ram_block3a581 = ram_block3a58_PORTADATAOUT_bus[0];

assign ram_block3a582 = ram_block3a58_PORTBDATAOUT_bus[0];

assign ram_block3a261 = ram_block3a26_PORTADATAOUT_bus[0];

assign ram_block3a262 = ram_block3a26_PORTBDATAOUT_bus[0];

assign ram_block3a591 = ram_block3a59_PORTADATAOUT_bus[0];

assign ram_block3a592 = ram_block3a59_PORTBDATAOUT_bus[0];

assign ram_block3a271 = ram_block3a27_PORTADATAOUT_bus[0];

assign ram_block3a272 = ram_block3a27_PORTBDATAOUT_bus[0];

assign ram_block3a601 = ram_block3a60_PORTADATAOUT_bus[0];

assign ram_block3a602 = ram_block3a60_PORTBDATAOUT_bus[0];

assign ram_block3a281 = ram_block3a28_PORTADATAOUT_bus[0];

assign ram_block3a282 = ram_block3a28_PORTBDATAOUT_bus[0];

assign ram_block3a611 = ram_block3a61_PORTADATAOUT_bus[0];

assign ram_block3a612 = ram_block3a61_PORTBDATAOUT_bus[0];

assign ram_block3a291 = ram_block3a29_PORTADATAOUT_bus[0];

assign ram_block3a292 = ram_block3a29_PORTBDATAOUT_bus[0];

assign ram_block3a621 = ram_block3a62_PORTADATAOUT_bus[0];

assign ram_block3a622 = ram_block3a62_PORTBDATAOUT_bus[0];

assign ram_block3a301 = ram_block3a30_PORTADATAOUT_bus[0];

assign ram_block3a302 = ram_block3a30_PORTBDATAOUT_bus[0];

assign ram_block3a631 = ram_block3a63_PORTADATAOUT_bus[0];

assign ram_block3a632 = ram_block3a63_PORTBDATAOUT_bus[0];

assign ram_block3a312 = ram_block3a31_PORTADATAOUT_bus[0];

assign ram_block3a313 = ram_block3a31_PORTBDATAOUT_bus[0];

decode_jsa_1 decode5(
	.ram_rom_addr_reg_13(ram_rom_addr_reg_13),
	.sdr(sdr),
	.eq_node_1(\decode5|eq_node[1]~0_combout ),
	.eq_node_0(\decode5|eq_node[0]~1_combout ),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

decode_jsa decode4(
	.ramaddr(ramaddr),
	.always1(always1),
	.ramWEN(ramWEN),
	.eq_node_1(\decode4|eq_node[1]~0_combout ),
	.eq_node_0(\decode4|eq_node[0]~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: M9K_X104_Y36_N0
cycloneive_ram_block ram_block3a32(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a32_PORTADATAOUT_bus),
	.portbdataout(ram_block3a32_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a32.clk0_core_clock_enable = "ena0";
defparam ram_block3a32.clk1_core_clock_enable = "ena1";
defparam ram_block3a32.data_interleave_offset_in_bits = 1;
defparam ram_block3a32.data_interleave_width_in_bits = 1;
defparam ram_block3a32.init_file = "meminit.hex";
defparam ram_block3a32.init_file_layout = "port_a";
defparam ram_block3a32.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a32.operation_mode = "bidir_dual_port";
defparam ram_block3a32.port_a_address_clear = "none";
defparam ram_block3a32.port_a_address_width = 13;
defparam ram_block3a32.port_a_byte_enable_clock = "none";
defparam ram_block3a32.port_a_data_out_clear = "none";
defparam ram_block3a32.port_a_data_out_clock = "none";
defparam ram_block3a32.port_a_data_width = 1;
defparam ram_block3a32.port_a_first_address = 0;
defparam ram_block3a32.port_a_first_bit_number = 0;
defparam ram_block3a32.port_a_last_address = 8191;
defparam ram_block3a32.port_a_logical_ram_depth = 16384;
defparam ram_block3a32.port_a_logical_ram_width = 32;
defparam ram_block3a32.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_address_clear = "none";
defparam ram_block3a32.port_b_address_clock = "clock1";
defparam ram_block3a32.port_b_address_width = 13;
defparam ram_block3a32.port_b_data_in_clock = "clock1";
defparam ram_block3a32.port_b_data_out_clear = "none";
defparam ram_block3a32.port_b_data_out_clock = "none";
defparam ram_block3a32.port_b_data_width = 1;
defparam ram_block3a32.port_b_first_address = 0;
defparam ram_block3a32.port_b_first_bit_number = 0;
defparam ram_block3a32.port_b_last_address = 8191;
defparam ram_block3a32.port_b_logical_ram_depth = 16384;
defparam ram_block3a32.port_b_logical_ram_width = 32;
defparam ram_block3a32.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_read_enable_clock = "clock1";
defparam ram_block3a32.port_b_write_enable_clock = "clock1";
defparam ram_block3a32.ram_block_type = "M9K";
defparam ram_block3a32.mem_init3 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007289B98206EA56527EF979635A0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y36_N0
cycloneive_ram_block ram_block3a0(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a0_PORTADATAOUT_bus),
	.portbdataout(ram_block3a0_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a0.clk0_core_clock_enable = "ena0";
defparam ram_block3a0.clk1_core_clock_enable = "ena1";
defparam ram_block3a0.data_interleave_offset_in_bits = 1;
defparam ram_block3a0.data_interleave_width_in_bits = 1;
defparam ram_block3a0.init_file = "meminit.hex";
defparam ram_block3a0.init_file_layout = "port_a";
defparam ram_block3a0.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a0.operation_mode = "bidir_dual_port";
defparam ram_block3a0.port_a_address_clear = "none";
defparam ram_block3a0.port_a_address_width = 13;
defparam ram_block3a0.port_a_byte_enable_clock = "none";
defparam ram_block3a0.port_a_data_out_clear = "none";
defparam ram_block3a0.port_a_data_out_clock = "none";
defparam ram_block3a0.port_a_data_width = 1;
defparam ram_block3a0.port_a_first_address = 0;
defparam ram_block3a0.port_a_first_bit_number = 0;
defparam ram_block3a0.port_a_last_address = 8191;
defparam ram_block3a0.port_a_logical_ram_depth = 16384;
defparam ram_block3a0.port_a_logical_ram_width = 32;
defparam ram_block3a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_address_clear = "none";
defparam ram_block3a0.port_b_address_clock = "clock1";
defparam ram_block3a0.port_b_address_width = 13;
defparam ram_block3a0.port_b_data_in_clock = "clock1";
defparam ram_block3a0.port_b_data_out_clear = "none";
defparam ram_block3a0.port_b_data_out_clock = "none";
defparam ram_block3a0.port_b_data_width = 1;
defparam ram_block3a0.port_b_first_address = 0;
defparam ram_block3a0.port_b_first_bit_number = 0;
defparam ram_block3a0.port_b_last_address = 8191;
defparam ram_block3a0.port_b_logical_ram_depth = 16384;
defparam ram_block3a0.port_b_logical_ram_width = 32;
defparam ram_block3a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_read_enable_clock = "clock1";
defparam ram_block3a0.port_b_write_enable_clock = "clock1";
defparam ram_block3a0.ram_block_type = "M9K";
defparam ram_block3a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011A02;
// synopsys translate_on

// Location: M9K_X104_Y41_N0
cycloneive_ram_block ram_block3a33(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a33_PORTADATAOUT_bus),
	.portbdataout(ram_block3a33_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a33.clk0_core_clock_enable = "ena0";
defparam ram_block3a33.clk1_core_clock_enable = "ena1";
defparam ram_block3a33.data_interleave_offset_in_bits = 1;
defparam ram_block3a33.data_interleave_width_in_bits = 1;
defparam ram_block3a33.init_file = "meminit.hex";
defparam ram_block3a33.init_file_layout = "port_a";
defparam ram_block3a33.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a33.operation_mode = "bidir_dual_port";
defparam ram_block3a33.port_a_address_clear = "none";
defparam ram_block3a33.port_a_address_width = 13;
defparam ram_block3a33.port_a_byte_enable_clock = "none";
defparam ram_block3a33.port_a_data_out_clear = "none";
defparam ram_block3a33.port_a_data_out_clock = "none";
defparam ram_block3a33.port_a_data_width = 1;
defparam ram_block3a33.port_a_first_address = 0;
defparam ram_block3a33.port_a_first_bit_number = 1;
defparam ram_block3a33.port_a_last_address = 8191;
defparam ram_block3a33.port_a_logical_ram_depth = 16384;
defparam ram_block3a33.port_a_logical_ram_width = 32;
defparam ram_block3a33.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_address_clear = "none";
defparam ram_block3a33.port_b_address_clock = "clock1";
defparam ram_block3a33.port_b_address_width = 13;
defparam ram_block3a33.port_b_data_in_clock = "clock1";
defparam ram_block3a33.port_b_data_out_clear = "none";
defparam ram_block3a33.port_b_data_out_clock = "none";
defparam ram_block3a33.port_b_data_width = 1;
defparam ram_block3a33.port_b_first_address = 0;
defparam ram_block3a33.port_b_first_bit_number = 1;
defparam ram_block3a33.port_b_last_address = 8191;
defparam ram_block3a33.port_b_logical_ram_depth = 16384;
defparam ram_block3a33.port_b_logical_ram_width = 32;
defparam ram_block3a33.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_read_enable_clock = "clock1";
defparam ram_block3a33.port_b_write_enable_clock = "clock1";
defparam ram_block3a33.ram_block_type = "M9K";
defparam ram_block3a33.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000592E61B5F6CACBDE18D9C2A9B20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X104_Y42_N0
cycloneive_ram_block ram_block3a1(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a1_PORTADATAOUT_bus),
	.portbdataout(ram_block3a1_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a1.clk0_core_clock_enable = "ena0";
defparam ram_block3a1.clk1_core_clock_enable = "ena1";
defparam ram_block3a1.data_interleave_offset_in_bits = 1;
defparam ram_block3a1.data_interleave_width_in_bits = 1;
defparam ram_block3a1.init_file = "meminit.hex";
defparam ram_block3a1.init_file_layout = "port_a";
defparam ram_block3a1.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a1.operation_mode = "bidir_dual_port";
defparam ram_block3a1.port_a_address_clear = "none";
defparam ram_block3a1.port_a_address_width = 13;
defparam ram_block3a1.port_a_byte_enable_clock = "none";
defparam ram_block3a1.port_a_data_out_clear = "none";
defparam ram_block3a1.port_a_data_out_clock = "none";
defparam ram_block3a1.port_a_data_width = 1;
defparam ram_block3a1.port_a_first_address = 0;
defparam ram_block3a1.port_a_first_bit_number = 1;
defparam ram_block3a1.port_a_last_address = 8191;
defparam ram_block3a1.port_a_logical_ram_depth = 16384;
defparam ram_block3a1.port_a_logical_ram_width = 32;
defparam ram_block3a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_address_clear = "none";
defparam ram_block3a1.port_b_address_clock = "clock1";
defparam ram_block3a1.port_b_address_width = 13;
defparam ram_block3a1.port_b_data_in_clock = "clock1";
defparam ram_block3a1.port_b_data_out_clear = "none";
defparam ram_block3a1.port_b_data_out_clock = "none";
defparam ram_block3a1.port_b_data_width = 1;
defparam ram_block3a1.port_b_first_address = 0;
defparam ram_block3a1.port_b_first_bit_number = 1;
defparam ram_block3a1.port_b_last_address = 8191;
defparam ram_block3a1.port_b_logical_ram_depth = 16384;
defparam ram_block3a1.port_b_logical_ram_width = 32;
defparam ram_block3a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_read_enable_clock = "clock1";
defparam ram_block3a1.port_b_write_enable_clock = "clock1";
defparam ram_block3a1.ram_block_type = "M9K";
defparam ram_block3a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013200;
// synopsys translate_on

// Location: M9K_X64_Y34_N0
cycloneive_ram_block ram_block3a34(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a34_PORTADATAOUT_bus),
	.portbdataout(ram_block3a34_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a34.clk0_core_clock_enable = "ena0";
defparam ram_block3a34.clk1_core_clock_enable = "ena1";
defparam ram_block3a34.data_interleave_offset_in_bits = 1;
defparam ram_block3a34.data_interleave_width_in_bits = 1;
defparam ram_block3a34.init_file = "meminit.hex";
defparam ram_block3a34.init_file_layout = "port_a";
defparam ram_block3a34.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a34.operation_mode = "bidir_dual_port";
defparam ram_block3a34.port_a_address_clear = "none";
defparam ram_block3a34.port_a_address_width = 13;
defparam ram_block3a34.port_a_byte_enable_clock = "none";
defparam ram_block3a34.port_a_data_out_clear = "none";
defparam ram_block3a34.port_a_data_out_clock = "none";
defparam ram_block3a34.port_a_data_width = 1;
defparam ram_block3a34.port_a_first_address = 0;
defparam ram_block3a34.port_a_first_bit_number = 2;
defparam ram_block3a34.port_a_last_address = 8191;
defparam ram_block3a34.port_a_logical_ram_depth = 16384;
defparam ram_block3a34.port_a_logical_ram_width = 32;
defparam ram_block3a34.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_address_clear = "none";
defparam ram_block3a34.port_b_address_clock = "clock1";
defparam ram_block3a34.port_b_address_width = 13;
defparam ram_block3a34.port_b_data_in_clock = "clock1";
defparam ram_block3a34.port_b_data_out_clear = "none";
defparam ram_block3a34.port_b_data_out_clock = "none";
defparam ram_block3a34.port_b_data_width = 1;
defparam ram_block3a34.port_b_first_address = 0;
defparam ram_block3a34.port_b_first_bit_number = 2;
defparam ram_block3a34.port_b_last_address = 8191;
defparam ram_block3a34.port_b_logical_ram_depth = 16384;
defparam ram_block3a34.port_b_logical_ram_width = 32;
defparam ram_block3a34.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_read_enable_clock = "clock1";
defparam ram_block3a34.port_b_write_enable_clock = "clock1";
defparam ram_block3a34.ram_block_type = "M9K";
defparam ram_block3a34.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000466F11FE97DE2DC7F80D940B0E0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y34_N0
cycloneive_ram_block ram_block3a2(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a2_PORTADATAOUT_bus),
	.portbdataout(ram_block3a2_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a2.clk0_core_clock_enable = "ena0";
defparam ram_block3a2.clk1_core_clock_enable = "ena1";
defparam ram_block3a2.data_interleave_offset_in_bits = 1;
defparam ram_block3a2.data_interleave_width_in_bits = 1;
defparam ram_block3a2.init_file = "meminit.hex";
defparam ram_block3a2.init_file_layout = "port_a";
defparam ram_block3a2.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a2.operation_mode = "bidir_dual_port";
defparam ram_block3a2.port_a_address_clear = "none";
defparam ram_block3a2.port_a_address_width = 13;
defparam ram_block3a2.port_a_byte_enable_clock = "none";
defparam ram_block3a2.port_a_data_out_clear = "none";
defparam ram_block3a2.port_a_data_out_clock = "none";
defparam ram_block3a2.port_a_data_width = 1;
defparam ram_block3a2.port_a_first_address = 0;
defparam ram_block3a2.port_a_first_bit_number = 2;
defparam ram_block3a2.port_a_last_address = 8191;
defparam ram_block3a2.port_a_logical_ram_depth = 16384;
defparam ram_block3a2.port_a_logical_ram_width = 32;
defparam ram_block3a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_address_clear = "none";
defparam ram_block3a2.port_b_address_clock = "clock1";
defparam ram_block3a2.port_b_address_width = 13;
defparam ram_block3a2.port_b_data_in_clock = "clock1";
defparam ram_block3a2.port_b_data_out_clear = "none";
defparam ram_block3a2.port_b_data_out_clock = "none";
defparam ram_block3a2.port_b_data_width = 1;
defparam ram_block3a2.port_b_first_address = 0;
defparam ram_block3a2.port_b_first_bit_number = 2;
defparam ram_block3a2.port_b_last_address = 8191;
defparam ram_block3a2.port_b_logical_ram_depth = 16384;
defparam ram_block3a2.port_b_logical_ram_width = 32;
defparam ram_block3a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_read_enable_clock = "clock1";
defparam ram_block3a2.port_b_write_enable_clock = "clock1";
defparam ram_block3a2.ram_block_type = "M9K";
defparam ram_block3a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010454;
// synopsys translate_on

// Location: M9K_X78_Y35_N0
cycloneive_ram_block ram_block3a35(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a35_PORTADATAOUT_bus),
	.portbdataout(ram_block3a35_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a35.clk0_core_clock_enable = "ena0";
defparam ram_block3a35.clk1_core_clock_enable = "ena1";
defparam ram_block3a35.data_interleave_offset_in_bits = 1;
defparam ram_block3a35.data_interleave_width_in_bits = 1;
defparam ram_block3a35.init_file = "meminit.hex";
defparam ram_block3a35.init_file_layout = "port_a";
defparam ram_block3a35.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a35.operation_mode = "bidir_dual_port";
defparam ram_block3a35.port_a_address_clear = "none";
defparam ram_block3a35.port_a_address_width = 13;
defparam ram_block3a35.port_a_byte_enable_clock = "none";
defparam ram_block3a35.port_a_data_out_clear = "none";
defparam ram_block3a35.port_a_data_out_clock = "none";
defparam ram_block3a35.port_a_data_width = 1;
defparam ram_block3a35.port_a_first_address = 0;
defparam ram_block3a35.port_a_first_bit_number = 3;
defparam ram_block3a35.port_a_last_address = 8191;
defparam ram_block3a35.port_a_logical_ram_depth = 16384;
defparam ram_block3a35.port_a_logical_ram_width = 32;
defparam ram_block3a35.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_address_clear = "none";
defparam ram_block3a35.port_b_address_clock = "clock1";
defparam ram_block3a35.port_b_address_width = 13;
defparam ram_block3a35.port_b_data_in_clock = "clock1";
defparam ram_block3a35.port_b_data_out_clear = "none";
defparam ram_block3a35.port_b_data_out_clock = "none";
defparam ram_block3a35.port_b_data_width = 1;
defparam ram_block3a35.port_b_first_address = 0;
defparam ram_block3a35.port_b_first_bit_number = 3;
defparam ram_block3a35.port_b_last_address = 8191;
defparam ram_block3a35.port_b_logical_ram_depth = 16384;
defparam ram_block3a35.port_b_logical_ram_width = 32;
defparam ram_block3a35.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_read_enable_clock = "clock1";
defparam ram_block3a35.port_b_write_enable_clock = "clock1";
defparam ram_block3a35.ram_block_type = "M9K";
defparam ram_block3a35.mem_init3 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000035B5D1D56E1A79B65BD7CACB7A0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y34_N0
cycloneive_ram_block ram_block3a3(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a3_PORTADATAOUT_bus),
	.portbdataout(ram_block3a3_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a3.clk0_core_clock_enable = "ena0";
defparam ram_block3a3.clk1_core_clock_enable = "ena1";
defparam ram_block3a3.data_interleave_offset_in_bits = 1;
defparam ram_block3a3.data_interleave_width_in_bits = 1;
defparam ram_block3a3.init_file = "meminit.hex";
defparam ram_block3a3.init_file_layout = "port_a";
defparam ram_block3a3.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a3.operation_mode = "bidir_dual_port";
defparam ram_block3a3.port_a_address_clear = "none";
defparam ram_block3a3.port_a_address_width = 13;
defparam ram_block3a3.port_a_byte_enable_clock = "none";
defparam ram_block3a3.port_a_data_out_clear = "none";
defparam ram_block3a3.port_a_data_out_clock = "none";
defparam ram_block3a3.port_a_data_width = 1;
defparam ram_block3a3.port_a_first_address = 0;
defparam ram_block3a3.port_a_first_bit_number = 3;
defparam ram_block3a3.port_a_last_address = 8191;
defparam ram_block3a3.port_a_logical_ram_depth = 16384;
defparam ram_block3a3.port_a_logical_ram_width = 32;
defparam ram_block3a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_address_clear = "none";
defparam ram_block3a3.port_b_address_clock = "clock1";
defparam ram_block3a3.port_b_address_width = 13;
defparam ram_block3a3.port_b_data_in_clock = "clock1";
defparam ram_block3a3.port_b_data_out_clear = "none";
defparam ram_block3a3.port_b_data_out_clock = "none";
defparam ram_block3a3.port_b_data_width = 1;
defparam ram_block3a3.port_b_first_address = 0;
defparam ram_block3a3.port_b_first_bit_number = 3;
defparam ram_block3a3.port_b_last_address = 8191;
defparam ram_block3a3.port_b_logical_ram_depth = 16384;
defparam ram_block3a3.port_b_logical_ram_width = 32;
defparam ram_block3a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_read_enable_clock = "clock1";
defparam ram_block3a3.port_b_write_enable_clock = "clock1";
defparam ram_block3a3.ram_block_type = "M9K";
defparam ram_block3a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014060;
// synopsys translate_on

// Location: M9K_X64_Y32_N0
cycloneive_ram_block ram_block3a36(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a36_PORTADATAOUT_bus),
	.portbdataout(ram_block3a36_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a36.clk0_core_clock_enable = "ena0";
defparam ram_block3a36.clk1_core_clock_enable = "ena1";
defparam ram_block3a36.data_interleave_offset_in_bits = 1;
defparam ram_block3a36.data_interleave_width_in_bits = 1;
defparam ram_block3a36.init_file = "meminit.hex";
defparam ram_block3a36.init_file_layout = "port_a";
defparam ram_block3a36.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a36.operation_mode = "bidir_dual_port";
defparam ram_block3a36.port_a_address_clear = "none";
defparam ram_block3a36.port_a_address_width = 13;
defparam ram_block3a36.port_a_byte_enable_clock = "none";
defparam ram_block3a36.port_a_data_out_clear = "none";
defparam ram_block3a36.port_a_data_out_clock = "none";
defparam ram_block3a36.port_a_data_width = 1;
defparam ram_block3a36.port_a_first_address = 0;
defparam ram_block3a36.port_a_first_bit_number = 4;
defparam ram_block3a36.port_a_last_address = 8191;
defparam ram_block3a36.port_a_logical_ram_depth = 16384;
defparam ram_block3a36.port_a_logical_ram_width = 32;
defparam ram_block3a36.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_address_clear = "none";
defparam ram_block3a36.port_b_address_clock = "clock1";
defparam ram_block3a36.port_b_address_width = 13;
defparam ram_block3a36.port_b_data_in_clock = "clock1";
defparam ram_block3a36.port_b_data_out_clear = "none";
defparam ram_block3a36.port_b_data_out_clock = "none";
defparam ram_block3a36.port_b_data_width = 1;
defparam ram_block3a36.port_b_first_address = 0;
defparam ram_block3a36.port_b_first_bit_number = 4;
defparam ram_block3a36.port_b_last_address = 8191;
defparam ram_block3a36.port_b_logical_ram_depth = 16384;
defparam ram_block3a36.port_b_logical_ram_width = 32;
defparam ram_block3a36.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_read_enable_clock = "clock1";
defparam ram_block3a36.port_b_write_enable_clock = "clock1";
defparam ram_block3a36.ram_block_type = "M9K";
defparam ram_block3a36.mem_init3 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000079A08B42BBB3DD751681DA88280000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y33_N0
cycloneive_ram_block ram_block3a4(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a4_PORTADATAOUT_bus),
	.portbdataout(ram_block3a4_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a4.clk0_core_clock_enable = "ena0";
defparam ram_block3a4.clk1_core_clock_enable = "ena1";
defparam ram_block3a4.data_interleave_offset_in_bits = 1;
defparam ram_block3a4.data_interleave_width_in_bits = 1;
defparam ram_block3a4.init_file = "meminit.hex";
defparam ram_block3a4.init_file_layout = "port_a";
defparam ram_block3a4.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a4.operation_mode = "bidir_dual_port";
defparam ram_block3a4.port_a_address_clear = "none";
defparam ram_block3a4.port_a_address_width = 13;
defparam ram_block3a4.port_a_byte_enable_clock = "none";
defparam ram_block3a4.port_a_data_out_clear = "none";
defparam ram_block3a4.port_a_data_out_clock = "none";
defparam ram_block3a4.port_a_data_width = 1;
defparam ram_block3a4.port_a_first_address = 0;
defparam ram_block3a4.port_a_first_bit_number = 4;
defparam ram_block3a4.port_a_last_address = 8191;
defparam ram_block3a4.port_a_logical_ram_depth = 16384;
defparam ram_block3a4.port_a_logical_ram_width = 32;
defparam ram_block3a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_address_clear = "none";
defparam ram_block3a4.port_b_address_clock = "clock1";
defparam ram_block3a4.port_b_address_width = 13;
defparam ram_block3a4.port_b_data_in_clock = "clock1";
defparam ram_block3a4.port_b_data_out_clear = "none";
defparam ram_block3a4.port_b_data_out_clock = "none";
defparam ram_block3a4.port_b_data_width = 1;
defparam ram_block3a4.port_b_first_address = 0;
defparam ram_block3a4.port_b_first_bit_number = 4;
defparam ram_block3a4.port_b_last_address = 8191;
defparam ram_block3a4.port_b_logical_ram_depth = 16384;
defparam ram_block3a4.port_b_logical_ram_width = 32;
defparam ram_block3a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_read_enable_clock = "clock1";
defparam ram_block3a4.port_b_write_enable_clock = "clock1";
defparam ram_block3a4.ram_block_type = "M9K";
defparam ram_block3a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014000;
// synopsys translate_on

// Location: M9K_X78_Y31_N0
cycloneive_ram_block ram_block3a37(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a37_PORTADATAOUT_bus),
	.portbdataout(ram_block3a37_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a37.clk0_core_clock_enable = "ena0";
defparam ram_block3a37.clk1_core_clock_enable = "ena1";
defparam ram_block3a37.data_interleave_offset_in_bits = 1;
defparam ram_block3a37.data_interleave_width_in_bits = 1;
defparam ram_block3a37.init_file = "meminit.hex";
defparam ram_block3a37.init_file_layout = "port_a";
defparam ram_block3a37.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a37.operation_mode = "bidir_dual_port";
defparam ram_block3a37.port_a_address_clear = "none";
defparam ram_block3a37.port_a_address_width = 13;
defparam ram_block3a37.port_a_byte_enable_clock = "none";
defparam ram_block3a37.port_a_data_out_clear = "none";
defparam ram_block3a37.port_a_data_out_clock = "none";
defparam ram_block3a37.port_a_data_width = 1;
defparam ram_block3a37.port_a_first_address = 0;
defparam ram_block3a37.port_a_first_bit_number = 5;
defparam ram_block3a37.port_a_last_address = 8191;
defparam ram_block3a37.port_a_logical_ram_depth = 16384;
defparam ram_block3a37.port_a_logical_ram_width = 32;
defparam ram_block3a37.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_address_clear = "none";
defparam ram_block3a37.port_b_address_clock = "clock1";
defparam ram_block3a37.port_b_address_width = 13;
defparam ram_block3a37.port_b_data_in_clock = "clock1";
defparam ram_block3a37.port_b_data_out_clear = "none";
defparam ram_block3a37.port_b_data_out_clock = "none";
defparam ram_block3a37.port_b_data_width = 1;
defparam ram_block3a37.port_b_first_address = 0;
defparam ram_block3a37.port_b_first_bit_number = 5;
defparam ram_block3a37.port_b_last_address = 8191;
defparam ram_block3a37.port_b_logical_ram_depth = 16384;
defparam ram_block3a37.port_b_logical_ram_width = 32;
defparam ram_block3a37.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_read_enable_clock = "clock1";
defparam ram_block3a37.port_b_write_enable_clock = "clock1";
defparam ram_block3a37.ram_block_type = "M9K";
defparam ram_block3a37.mem_init3 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006A801AC0C797222BAD3D00668E0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y33_N0
cycloneive_ram_block ram_block3a5(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a5_PORTADATAOUT_bus),
	.portbdataout(ram_block3a5_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a5.clk0_core_clock_enable = "ena0";
defparam ram_block3a5.clk1_core_clock_enable = "ena1";
defparam ram_block3a5.data_interleave_offset_in_bits = 1;
defparam ram_block3a5.data_interleave_width_in_bits = 1;
defparam ram_block3a5.init_file = "meminit.hex";
defparam ram_block3a5.init_file_layout = "port_a";
defparam ram_block3a5.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a5.operation_mode = "bidir_dual_port";
defparam ram_block3a5.port_a_address_clear = "none";
defparam ram_block3a5.port_a_address_width = 13;
defparam ram_block3a5.port_a_byte_enable_clock = "none";
defparam ram_block3a5.port_a_data_out_clear = "none";
defparam ram_block3a5.port_a_data_out_clock = "none";
defparam ram_block3a5.port_a_data_width = 1;
defparam ram_block3a5.port_a_first_address = 0;
defparam ram_block3a5.port_a_first_bit_number = 5;
defparam ram_block3a5.port_a_last_address = 8191;
defparam ram_block3a5.port_a_logical_ram_depth = 16384;
defparam ram_block3a5.port_a_logical_ram_width = 32;
defparam ram_block3a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_address_clear = "none";
defparam ram_block3a5.port_b_address_clock = "clock1";
defparam ram_block3a5.port_b_address_width = 13;
defparam ram_block3a5.port_b_data_in_clock = "clock1";
defparam ram_block3a5.port_b_data_out_clear = "none";
defparam ram_block3a5.port_b_data_out_clock = "none";
defparam ram_block3a5.port_b_data_width = 1;
defparam ram_block3a5.port_b_first_address = 0;
defparam ram_block3a5.port_b_first_bit_number = 5;
defparam ram_block3a5.port_b_last_address = 8191;
defparam ram_block3a5.port_b_logical_ram_depth = 16384;
defparam ram_block3a5.port_b_logical_ram_width = 32;
defparam ram_block3a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_read_enable_clock = "clock1";
defparam ram_block3a5.port_b_write_enable_clock = "clock1";
defparam ram_block3a5.ram_block_type = "M9K";
defparam ram_block3a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000015A00;
// synopsys translate_on

// Location: M9K_X64_Y41_N0
cycloneive_ram_block ram_block3a38(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a38_PORTADATAOUT_bus),
	.portbdataout(ram_block3a38_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a38.clk0_core_clock_enable = "ena0";
defparam ram_block3a38.clk1_core_clock_enable = "ena1";
defparam ram_block3a38.data_interleave_offset_in_bits = 1;
defparam ram_block3a38.data_interleave_width_in_bits = 1;
defparam ram_block3a38.init_file = "meminit.hex";
defparam ram_block3a38.init_file_layout = "port_a";
defparam ram_block3a38.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a38.operation_mode = "bidir_dual_port";
defparam ram_block3a38.port_a_address_clear = "none";
defparam ram_block3a38.port_a_address_width = 13;
defparam ram_block3a38.port_a_byte_enable_clock = "none";
defparam ram_block3a38.port_a_data_out_clear = "none";
defparam ram_block3a38.port_a_data_out_clock = "none";
defparam ram_block3a38.port_a_data_width = 1;
defparam ram_block3a38.port_a_first_address = 0;
defparam ram_block3a38.port_a_first_bit_number = 6;
defparam ram_block3a38.port_a_last_address = 8191;
defparam ram_block3a38.port_a_logical_ram_depth = 16384;
defparam ram_block3a38.port_a_logical_ram_width = 32;
defparam ram_block3a38.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_address_clear = "none";
defparam ram_block3a38.port_b_address_clock = "clock1";
defparam ram_block3a38.port_b_address_width = 13;
defparam ram_block3a38.port_b_data_in_clock = "clock1";
defparam ram_block3a38.port_b_data_out_clear = "none";
defparam ram_block3a38.port_b_data_out_clock = "none";
defparam ram_block3a38.port_b_data_width = 1;
defparam ram_block3a38.port_b_first_address = 0;
defparam ram_block3a38.port_b_first_bit_number = 6;
defparam ram_block3a38.port_b_last_address = 8191;
defparam ram_block3a38.port_b_logical_ram_depth = 16384;
defparam ram_block3a38.port_b_logical_ram_width = 32;
defparam ram_block3a38.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_read_enable_clock = "clock1";
defparam ram_block3a38.port_b_write_enable_clock = "clock1";
defparam ram_block3a38.ram_block_type = "M9K";
defparam ram_block3a38.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000711CAD5E440ED8933DD8400E1E0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y44_N0
cycloneive_ram_block ram_block3a6(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a6_PORTADATAOUT_bus),
	.portbdataout(ram_block3a6_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a6.clk0_core_clock_enable = "ena0";
defparam ram_block3a6.clk1_core_clock_enable = "ena1";
defparam ram_block3a6.data_interleave_offset_in_bits = 1;
defparam ram_block3a6.data_interleave_width_in_bits = 1;
defparam ram_block3a6.init_file = "meminit.hex";
defparam ram_block3a6.init_file_layout = "port_a";
defparam ram_block3a6.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a6.operation_mode = "bidir_dual_port";
defparam ram_block3a6.port_a_address_clear = "none";
defparam ram_block3a6.port_a_address_width = 13;
defparam ram_block3a6.port_a_byte_enable_clock = "none";
defparam ram_block3a6.port_a_data_out_clear = "none";
defparam ram_block3a6.port_a_data_out_clock = "none";
defparam ram_block3a6.port_a_data_width = 1;
defparam ram_block3a6.port_a_first_address = 0;
defparam ram_block3a6.port_a_first_bit_number = 6;
defparam ram_block3a6.port_a_last_address = 8191;
defparam ram_block3a6.port_a_logical_ram_depth = 16384;
defparam ram_block3a6.port_a_logical_ram_width = 32;
defparam ram_block3a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_address_clear = "none";
defparam ram_block3a6.port_b_address_clock = "clock1";
defparam ram_block3a6.port_b_address_width = 13;
defparam ram_block3a6.port_b_data_in_clock = "clock1";
defparam ram_block3a6.port_b_data_out_clear = "none";
defparam ram_block3a6.port_b_data_out_clock = "none";
defparam ram_block3a6.port_b_data_width = 1;
defparam ram_block3a6.port_b_first_address = 0;
defparam ram_block3a6.port_b_first_bit_number = 6;
defparam ram_block3a6.port_b_last_address = 8191;
defparam ram_block3a6.port_b_logical_ram_depth = 16384;
defparam ram_block3a6.port_b_logical_ram_width = 32;
defparam ram_block3a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_read_enable_clock = "clock1";
defparam ram_block3a6.port_b_write_enable_clock = "clock1";
defparam ram_block3a6.ram_block_type = "M9K";
defparam ram_block3a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014000;
// synopsys translate_on

// Location: M9K_X104_Y39_N0
cycloneive_ram_block ram_block3a39(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a39_PORTADATAOUT_bus),
	.portbdataout(ram_block3a39_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a39.clk0_core_clock_enable = "ena0";
defparam ram_block3a39.clk1_core_clock_enable = "ena1";
defparam ram_block3a39.data_interleave_offset_in_bits = 1;
defparam ram_block3a39.data_interleave_width_in_bits = 1;
defparam ram_block3a39.init_file = "meminit.hex";
defparam ram_block3a39.init_file_layout = "port_a";
defparam ram_block3a39.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a39.operation_mode = "bidir_dual_port";
defparam ram_block3a39.port_a_address_clear = "none";
defparam ram_block3a39.port_a_address_width = 13;
defparam ram_block3a39.port_a_byte_enable_clock = "none";
defparam ram_block3a39.port_a_data_out_clear = "none";
defparam ram_block3a39.port_a_data_out_clock = "none";
defparam ram_block3a39.port_a_data_width = 1;
defparam ram_block3a39.port_a_first_address = 0;
defparam ram_block3a39.port_a_first_bit_number = 7;
defparam ram_block3a39.port_a_last_address = 8191;
defparam ram_block3a39.port_a_logical_ram_depth = 16384;
defparam ram_block3a39.port_a_logical_ram_width = 32;
defparam ram_block3a39.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_address_clear = "none";
defparam ram_block3a39.port_b_address_clock = "clock1";
defparam ram_block3a39.port_b_address_width = 13;
defparam ram_block3a39.port_b_data_in_clock = "clock1";
defparam ram_block3a39.port_b_data_out_clear = "none";
defparam ram_block3a39.port_b_data_out_clock = "none";
defparam ram_block3a39.port_b_data_width = 1;
defparam ram_block3a39.port_b_first_address = 0;
defparam ram_block3a39.port_b_first_bit_number = 7;
defparam ram_block3a39.port_b_last_address = 8191;
defparam ram_block3a39.port_b_logical_ram_depth = 16384;
defparam ram_block3a39.port_b_logical_ram_width = 32;
defparam ram_block3a39.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_read_enable_clock = "clock1";
defparam ram_block3a39.port_b_write_enable_clock = "clock1";
defparam ram_block3a39.ram_block_type = "M9K";
defparam ram_block3a39.mem_init3 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000078E4785C3A8D6790D22EAF70100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y39_N0
cycloneive_ram_block ram_block3a7(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a7_PORTADATAOUT_bus),
	.portbdataout(ram_block3a7_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a7.clk0_core_clock_enable = "ena0";
defparam ram_block3a7.clk1_core_clock_enable = "ena1";
defparam ram_block3a7.data_interleave_offset_in_bits = 1;
defparam ram_block3a7.data_interleave_width_in_bits = 1;
defparam ram_block3a7.init_file = "meminit.hex";
defparam ram_block3a7.init_file_layout = "port_a";
defparam ram_block3a7.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a7.operation_mode = "bidir_dual_port";
defparam ram_block3a7.port_a_address_clear = "none";
defparam ram_block3a7.port_a_address_width = 13;
defparam ram_block3a7.port_a_byte_enable_clock = "none";
defparam ram_block3a7.port_a_data_out_clear = "none";
defparam ram_block3a7.port_a_data_out_clock = "none";
defparam ram_block3a7.port_a_data_width = 1;
defparam ram_block3a7.port_a_first_address = 0;
defparam ram_block3a7.port_a_first_bit_number = 7;
defparam ram_block3a7.port_a_last_address = 8191;
defparam ram_block3a7.port_a_logical_ram_depth = 16384;
defparam ram_block3a7.port_a_logical_ram_width = 32;
defparam ram_block3a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_address_clear = "none";
defparam ram_block3a7.port_b_address_clock = "clock1";
defparam ram_block3a7.port_b_address_width = 13;
defparam ram_block3a7.port_b_data_in_clock = "clock1";
defparam ram_block3a7.port_b_data_out_clear = "none";
defparam ram_block3a7.port_b_data_out_clock = "none";
defparam ram_block3a7.port_b_data_width = 1;
defparam ram_block3a7.port_b_first_address = 0;
defparam ram_block3a7.port_b_first_bit_number = 7;
defparam ram_block3a7.port_b_last_address = 8191;
defparam ram_block3a7.port_b_logical_ram_depth = 16384;
defparam ram_block3a7.port_b_logical_ram_width = 32;
defparam ram_block3a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_read_enable_clock = "clock1";
defparam ram_block3a7.port_b_write_enable_clock = "clock1";
defparam ram_block3a7.ram_block_type = "M9K";
defparam ram_block3a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014000;
// synopsys translate_on

// Location: M9K_X104_Y40_N0
cycloneive_ram_block ram_block3a40(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a40_PORTADATAOUT_bus),
	.portbdataout(ram_block3a40_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a40.clk0_core_clock_enable = "ena0";
defparam ram_block3a40.clk1_core_clock_enable = "ena1";
defparam ram_block3a40.data_interleave_offset_in_bits = 1;
defparam ram_block3a40.data_interleave_width_in_bits = 1;
defparam ram_block3a40.init_file = "meminit.hex";
defparam ram_block3a40.init_file_layout = "port_a";
defparam ram_block3a40.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a40.operation_mode = "bidir_dual_port";
defparam ram_block3a40.port_a_address_clear = "none";
defparam ram_block3a40.port_a_address_width = 13;
defparam ram_block3a40.port_a_byte_enable_clock = "none";
defparam ram_block3a40.port_a_data_out_clear = "none";
defparam ram_block3a40.port_a_data_out_clock = "none";
defparam ram_block3a40.port_a_data_width = 1;
defparam ram_block3a40.port_a_first_address = 0;
defparam ram_block3a40.port_a_first_bit_number = 8;
defparam ram_block3a40.port_a_last_address = 8191;
defparam ram_block3a40.port_a_logical_ram_depth = 16384;
defparam ram_block3a40.port_a_logical_ram_width = 32;
defparam ram_block3a40.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_address_clear = "none";
defparam ram_block3a40.port_b_address_clock = "clock1";
defparam ram_block3a40.port_b_address_width = 13;
defparam ram_block3a40.port_b_data_in_clock = "clock1";
defparam ram_block3a40.port_b_data_out_clear = "none";
defparam ram_block3a40.port_b_data_out_clock = "none";
defparam ram_block3a40.port_b_data_width = 1;
defparam ram_block3a40.port_b_first_address = 0;
defparam ram_block3a40.port_b_first_bit_number = 8;
defparam ram_block3a40.port_b_last_address = 8191;
defparam ram_block3a40.port_b_logical_ram_depth = 16384;
defparam ram_block3a40.port_b_logical_ram_width = 32;
defparam ram_block3a40.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_read_enable_clock = "clock1";
defparam ram_block3a40.port_b_write_enable_clock = "clock1";
defparam ram_block3a40.ram_block_type = "M9K";
defparam ram_block3a40.mem_init3 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000024B0BEB5CD48A0C4A466CF94D00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X104_Y37_N0
cycloneive_ram_block ram_block3a8(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a8_PORTADATAOUT_bus),
	.portbdataout(ram_block3a8_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a8.clk0_core_clock_enable = "ena0";
defparam ram_block3a8.clk1_core_clock_enable = "ena1";
defparam ram_block3a8.data_interleave_offset_in_bits = 1;
defparam ram_block3a8.data_interleave_width_in_bits = 1;
defparam ram_block3a8.init_file = "meminit.hex";
defparam ram_block3a8.init_file_layout = "port_a";
defparam ram_block3a8.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a8.operation_mode = "bidir_dual_port";
defparam ram_block3a8.port_a_address_clear = "none";
defparam ram_block3a8.port_a_address_width = 13;
defparam ram_block3a8.port_a_byte_enable_clock = "none";
defparam ram_block3a8.port_a_data_out_clear = "none";
defparam ram_block3a8.port_a_data_out_clock = "none";
defparam ram_block3a8.port_a_data_width = 1;
defparam ram_block3a8.port_a_first_address = 0;
defparam ram_block3a8.port_a_first_bit_number = 8;
defparam ram_block3a8.port_a_last_address = 8191;
defparam ram_block3a8.port_a_logical_ram_depth = 16384;
defparam ram_block3a8.port_a_logical_ram_width = 32;
defparam ram_block3a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_address_clear = "none";
defparam ram_block3a8.port_b_address_clock = "clock1";
defparam ram_block3a8.port_b_address_width = 13;
defparam ram_block3a8.port_b_data_in_clock = "clock1";
defparam ram_block3a8.port_b_data_out_clear = "none";
defparam ram_block3a8.port_b_data_out_clock = "none";
defparam ram_block3a8.port_b_data_width = 1;
defparam ram_block3a8.port_b_first_address = 0;
defparam ram_block3a8.port_b_first_bit_number = 8;
defparam ram_block3a8.port_b_last_address = 8191;
defparam ram_block3a8.port_b_logical_ram_depth = 16384;
defparam ram_block3a8.port_b_logical_ram_width = 32;
defparam ram_block3a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_read_enable_clock = "clock1";
defparam ram_block3a8.port_b_write_enable_clock = "clock1";
defparam ram_block3a8.ram_block_type = "M9K";
defparam ram_block3a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014000;
// synopsys translate_on

// Location: M9K_X64_Y40_N0
cycloneive_ram_block ram_block3a41(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a41_PORTADATAOUT_bus),
	.portbdataout(ram_block3a41_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a41.clk0_core_clock_enable = "ena0";
defparam ram_block3a41.clk1_core_clock_enable = "ena1";
defparam ram_block3a41.data_interleave_offset_in_bits = 1;
defparam ram_block3a41.data_interleave_width_in_bits = 1;
defparam ram_block3a41.init_file = "meminit.hex";
defparam ram_block3a41.init_file_layout = "port_a";
defparam ram_block3a41.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a41.operation_mode = "bidir_dual_port";
defparam ram_block3a41.port_a_address_clear = "none";
defparam ram_block3a41.port_a_address_width = 13;
defparam ram_block3a41.port_a_byte_enable_clock = "none";
defparam ram_block3a41.port_a_data_out_clear = "none";
defparam ram_block3a41.port_a_data_out_clock = "none";
defparam ram_block3a41.port_a_data_width = 1;
defparam ram_block3a41.port_a_first_address = 0;
defparam ram_block3a41.port_a_first_bit_number = 9;
defparam ram_block3a41.port_a_last_address = 8191;
defparam ram_block3a41.port_a_logical_ram_depth = 16384;
defparam ram_block3a41.port_a_logical_ram_width = 32;
defparam ram_block3a41.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_address_clear = "none";
defparam ram_block3a41.port_b_address_clock = "clock1";
defparam ram_block3a41.port_b_address_width = 13;
defparam ram_block3a41.port_b_data_in_clock = "clock1";
defparam ram_block3a41.port_b_data_out_clear = "none";
defparam ram_block3a41.port_b_data_out_clock = "none";
defparam ram_block3a41.port_b_data_width = 1;
defparam ram_block3a41.port_b_first_address = 0;
defparam ram_block3a41.port_b_first_bit_number = 9;
defparam ram_block3a41.port_b_last_address = 8191;
defparam ram_block3a41.port_b_logical_ram_depth = 16384;
defparam ram_block3a41.port_b_logical_ram_width = 32;
defparam ram_block3a41.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_read_enable_clock = "clock1";
defparam ram_block3a41.port_b_write_enable_clock = "clock1";
defparam ram_block3a41.ram_block_type = "M9K";
defparam ram_block3a41.mem_init3 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006E16818E27D32BC984B5234E100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y40_N0
cycloneive_ram_block ram_block3a9(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a9_PORTADATAOUT_bus),
	.portbdataout(ram_block3a9_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a9.clk0_core_clock_enable = "ena0";
defparam ram_block3a9.clk1_core_clock_enable = "ena1";
defparam ram_block3a9.data_interleave_offset_in_bits = 1;
defparam ram_block3a9.data_interleave_width_in_bits = 1;
defparam ram_block3a9.init_file = "meminit.hex";
defparam ram_block3a9.init_file_layout = "port_a";
defparam ram_block3a9.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a9.operation_mode = "bidir_dual_port";
defparam ram_block3a9.port_a_address_clear = "none";
defparam ram_block3a9.port_a_address_width = 13;
defparam ram_block3a9.port_a_byte_enable_clock = "none";
defparam ram_block3a9.port_a_data_out_clear = "none";
defparam ram_block3a9.port_a_data_out_clock = "none";
defparam ram_block3a9.port_a_data_width = 1;
defparam ram_block3a9.port_a_first_address = 0;
defparam ram_block3a9.port_a_first_bit_number = 9;
defparam ram_block3a9.port_a_last_address = 8191;
defparam ram_block3a9.port_a_logical_ram_depth = 16384;
defparam ram_block3a9.port_a_logical_ram_width = 32;
defparam ram_block3a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_address_clear = "none";
defparam ram_block3a9.port_b_address_clock = "clock1";
defparam ram_block3a9.port_b_address_width = 13;
defparam ram_block3a9.port_b_data_in_clock = "clock1";
defparam ram_block3a9.port_b_data_out_clear = "none";
defparam ram_block3a9.port_b_data_out_clock = "none";
defparam ram_block3a9.port_b_data_width = 1;
defparam ram_block3a9.port_b_first_address = 0;
defparam ram_block3a9.port_b_first_bit_number = 9;
defparam ram_block3a9.port_b_last_address = 8191;
defparam ram_block3a9.port_b_logical_ram_depth = 16384;
defparam ram_block3a9.port_b_logical_ram_width = 32;
defparam ram_block3a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_read_enable_clock = "clock1";
defparam ram_block3a9.port_b_write_enable_clock = "clock1";
defparam ram_block3a9.ram_block_type = "M9K";
defparam ram_block3a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014000;
// synopsys translate_on

// Location: M9K_X78_Y37_N0
cycloneive_ram_block ram_block3a42(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a42_PORTADATAOUT_bus),
	.portbdataout(ram_block3a42_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a42.clk0_core_clock_enable = "ena0";
defparam ram_block3a42.clk1_core_clock_enable = "ena1";
defparam ram_block3a42.data_interleave_offset_in_bits = 1;
defparam ram_block3a42.data_interleave_width_in_bits = 1;
defparam ram_block3a42.init_file = "meminit.hex";
defparam ram_block3a42.init_file_layout = "port_a";
defparam ram_block3a42.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a42.operation_mode = "bidir_dual_port";
defparam ram_block3a42.port_a_address_clear = "none";
defparam ram_block3a42.port_a_address_width = 13;
defparam ram_block3a42.port_a_byte_enable_clock = "none";
defparam ram_block3a42.port_a_data_out_clear = "none";
defparam ram_block3a42.port_a_data_out_clock = "none";
defparam ram_block3a42.port_a_data_width = 1;
defparam ram_block3a42.port_a_first_address = 0;
defparam ram_block3a42.port_a_first_bit_number = 10;
defparam ram_block3a42.port_a_last_address = 8191;
defparam ram_block3a42.port_a_logical_ram_depth = 16384;
defparam ram_block3a42.port_a_logical_ram_width = 32;
defparam ram_block3a42.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_address_clear = "none";
defparam ram_block3a42.port_b_address_clock = "clock1";
defparam ram_block3a42.port_b_address_width = 13;
defparam ram_block3a42.port_b_data_in_clock = "clock1";
defparam ram_block3a42.port_b_data_out_clear = "none";
defparam ram_block3a42.port_b_data_out_clock = "none";
defparam ram_block3a42.port_b_data_width = 1;
defparam ram_block3a42.port_b_first_address = 0;
defparam ram_block3a42.port_b_first_bit_number = 10;
defparam ram_block3a42.port_b_last_address = 8191;
defparam ram_block3a42.port_b_logical_ram_depth = 16384;
defparam ram_block3a42.port_b_logical_ram_width = 32;
defparam ram_block3a42.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_read_enable_clock = "clock1";
defparam ram_block3a42.port_b_write_enable_clock = "clock1";
defparam ram_block3a42.ram_block_type = "M9K";
defparam ram_block3a42.mem_init3 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010993F705D79849316AA6F56B20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X104_Y38_N0
cycloneive_ram_block ram_block3a10(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a10_PORTADATAOUT_bus),
	.portbdataout(ram_block3a10_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a10.clk0_core_clock_enable = "ena0";
defparam ram_block3a10.clk1_core_clock_enable = "ena1";
defparam ram_block3a10.data_interleave_offset_in_bits = 1;
defparam ram_block3a10.data_interleave_width_in_bits = 1;
defparam ram_block3a10.init_file = "meminit.hex";
defparam ram_block3a10.init_file_layout = "port_a";
defparam ram_block3a10.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a10.operation_mode = "bidir_dual_port";
defparam ram_block3a10.port_a_address_clear = "none";
defparam ram_block3a10.port_a_address_width = 13;
defparam ram_block3a10.port_a_byte_enable_clock = "none";
defparam ram_block3a10.port_a_data_out_clear = "none";
defparam ram_block3a10.port_a_data_out_clock = "none";
defparam ram_block3a10.port_a_data_width = 1;
defparam ram_block3a10.port_a_first_address = 0;
defparam ram_block3a10.port_a_first_bit_number = 10;
defparam ram_block3a10.port_a_last_address = 8191;
defparam ram_block3a10.port_a_logical_ram_depth = 16384;
defparam ram_block3a10.port_a_logical_ram_width = 32;
defparam ram_block3a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_address_clear = "none";
defparam ram_block3a10.port_b_address_clock = "clock1";
defparam ram_block3a10.port_b_address_width = 13;
defparam ram_block3a10.port_b_data_in_clock = "clock1";
defparam ram_block3a10.port_b_data_out_clear = "none";
defparam ram_block3a10.port_b_data_out_clock = "none";
defparam ram_block3a10.port_b_data_width = 1;
defparam ram_block3a10.port_b_first_address = 0;
defparam ram_block3a10.port_b_first_bit_number = 10;
defparam ram_block3a10.port_b_last_address = 8191;
defparam ram_block3a10.port_b_logical_ram_depth = 16384;
defparam ram_block3a10.port_b_logical_ram_width = 32;
defparam ram_block3a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_read_enable_clock = "clock1";
defparam ram_block3a10.port_b_write_enable_clock = "clock1";
defparam ram_block3a10.ram_block_type = "M9K";
defparam ram_block3a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014000;
// synopsys translate_on

// Location: M9K_X64_Y39_N0
cycloneive_ram_block ram_block3a43(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a43_PORTADATAOUT_bus),
	.portbdataout(ram_block3a43_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a43.clk0_core_clock_enable = "ena0";
defparam ram_block3a43.clk1_core_clock_enable = "ena1";
defparam ram_block3a43.data_interleave_offset_in_bits = 1;
defparam ram_block3a43.data_interleave_width_in_bits = 1;
defparam ram_block3a43.init_file = "meminit.hex";
defparam ram_block3a43.init_file_layout = "port_a";
defparam ram_block3a43.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a43.operation_mode = "bidir_dual_port";
defparam ram_block3a43.port_a_address_clear = "none";
defparam ram_block3a43.port_a_address_width = 13;
defparam ram_block3a43.port_a_byte_enable_clock = "none";
defparam ram_block3a43.port_a_data_out_clear = "none";
defparam ram_block3a43.port_a_data_out_clock = "none";
defparam ram_block3a43.port_a_data_width = 1;
defparam ram_block3a43.port_a_first_address = 0;
defparam ram_block3a43.port_a_first_bit_number = 11;
defparam ram_block3a43.port_a_last_address = 8191;
defparam ram_block3a43.port_a_logical_ram_depth = 16384;
defparam ram_block3a43.port_a_logical_ram_width = 32;
defparam ram_block3a43.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_address_clear = "none";
defparam ram_block3a43.port_b_address_clock = "clock1";
defparam ram_block3a43.port_b_address_width = 13;
defparam ram_block3a43.port_b_data_in_clock = "clock1";
defparam ram_block3a43.port_b_data_out_clear = "none";
defparam ram_block3a43.port_b_data_out_clock = "none";
defparam ram_block3a43.port_b_data_width = 1;
defparam ram_block3a43.port_b_first_address = 0;
defparam ram_block3a43.port_b_first_bit_number = 11;
defparam ram_block3a43.port_b_last_address = 8191;
defparam ram_block3a43.port_b_logical_ram_depth = 16384;
defparam ram_block3a43.port_b_logical_ram_width = 32;
defparam ram_block3a43.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_read_enable_clock = "clock1";
defparam ram_block3a43.port_b_write_enable_clock = "clock1";
defparam ram_block3a43.ram_block_type = "M9K";
defparam ram_block3a43.mem_init3 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000024B613BE67C43B53C478A34C1A0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y43_N0
cycloneive_ram_block ram_block3a11(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a11_PORTADATAOUT_bus),
	.portbdataout(ram_block3a11_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a11.clk0_core_clock_enable = "ena0";
defparam ram_block3a11.clk1_core_clock_enable = "ena1";
defparam ram_block3a11.data_interleave_offset_in_bits = 1;
defparam ram_block3a11.data_interleave_width_in_bits = 1;
defparam ram_block3a11.init_file = "meminit.hex";
defparam ram_block3a11.init_file_layout = "port_a";
defparam ram_block3a11.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a11.operation_mode = "bidir_dual_port";
defparam ram_block3a11.port_a_address_clear = "none";
defparam ram_block3a11.port_a_address_width = 13;
defparam ram_block3a11.port_a_byte_enable_clock = "none";
defparam ram_block3a11.port_a_data_out_clear = "none";
defparam ram_block3a11.port_a_data_out_clock = "none";
defparam ram_block3a11.port_a_data_width = 1;
defparam ram_block3a11.port_a_first_address = 0;
defparam ram_block3a11.port_a_first_bit_number = 11;
defparam ram_block3a11.port_a_last_address = 8191;
defparam ram_block3a11.port_a_logical_ram_depth = 16384;
defparam ram_block3a11.port_a_logical_ram_width = 32;
defparam ram_block3a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_address_clear = "none";
defparam ram_block3a11.port_b_address_clock = "clock1";
defparam ram_block3a11.port_b_address_width = 13;
defparam ram_block3a11.port_b_data_in_clock = "clock1";
defparam ram_block3a11.port_b_data_out_clear = "none";
defparam ram_block3a11.port_b_data_out_clock = "none";
defparam ram_block3a11.port_b_data_width = 1;
defparam ram_block3a11.port_b_first_address = 0;
defparam ram_block3a11.port_b_first_bit_number = 11;
defparam ram_block3a11.port_b_last_address = 8191;
defparam ram_block3a11.port_b_logical_ram_depth = 16384;
defparam ram_block3a11.port_b_logical_ram_width = 32;
defparam ram_block3a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_read_enable_clock = "clock1";
defparam ram_block3a11.port_b_write_enable_clock = "clock1";
defparam ram_block3a11.ram_block_type = "M9K";
defparam ram_block3a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014A00;
// synopsys translate_on

// Location: M9K_X104_Y43_N0
cycloneive_ram_block ram_block3a44(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a44_PORTADATAOUT_bus),
	.portbdataout(ram_block3a44_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a44.clk0_core_clock_enable = "ena0";
defparam ram_block3a44.clk1_core_clock_enable = "ena1";
defparam ram_block3a44.data_interleave_offset_in_bits = 1;
defparam ram_block3a44.data_interleave_width_in_bits = 1;
defparam ram_block3a44.init_file = "meminit.hex";
defparam ram_block3a44.init_file_layout = "port_a";
defparam ram_block3a44.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a44.operation_mode = "bidir_dual_port";
defparam ram_block3a44.port_a_address_clear = "none";
defparam ram_block3a44.port_a_address_width = 13;
defparam ram_block3a44.port_a_byte_enable_clock = "none";
defparam ram_block3a44.port_a_data_out_clear = "none";
defparam ram_block3a44.port_a_data_out_clock = "none";
defparam ram_block3a44.port_a_data_width = 1;
defparam ram_block3a44.port_a_first_address = 0;
defparam ram_block3a44.port_a_first_bit_number = 12;
defparam ram_block3a44.port_a_last_address = 8191;
defparam ram_block3a44.port_a_logical_ram_depth = 16384;
defparam ram_block3a44.port_a_logical_ram_width = 32;
defparam ram_block3a44.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_address_clear = "none";
defparam ram_block3a44.port_b_address_clock = "clock1";
defparam ram_block3a44.port_b_address_width = 13;
defparam ram_block3a44.port_b_data_in_clock = "clock1";
defparam ram_block3a44.port_b_data_out_clear = "none";
defparam ram_block3a44.port_b_data_out_clock = "none";
defparam ram_block3a44.port_b_data_width = 1;
defparam ram_block3a44.port_b_first_address = 0;
defparam ram_block3a44.port_b_first_bit_number = 12;
defparam ram_block3a44.port_b_last_address = 8191;
defparam ram_block3a44.port_b_logical_ram_depth = 16384;
defparam ram_block3a44.port_b_logical_ram_width = 32;
defparam ram_block3a44.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_read_enable_clock = "clock1";
defparam ram_block3a44.port_b_write_enable_clock = "clock1";
defparam ram_block3a44.ram_block_type = "M9K";
defparam ram_block3a44.mem_init3 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004C9F5AB072B2D6AE7E2EC0B3120000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y39_N0
cycloneive_ram_block ram_block3a12(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a12_PORTADATAOUT_bus),
	.portbdataout(ram_block3a12_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a12.clk0_core_clock_enable = "ena0";
defparam ram_block3a12.clk1_core_clock_enable = "ena1";
defparam ram_block3a12.data_interleave_offset_in_bits = 1;
defparam ram_block3a12.data_interleave_width_in_bits = 1;
defparam ram_block3a12.init_file = "meminit.hex";
defparam ram_block3a12.init_file_layout = "port_a";
defparam ram_block3a12.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a12.operation_mode = "bidir_dual_port";
defparam ram_block3a12.port_a_address_clear = "none";
defparam ram_block3a12.port_a_address_width = 13;
defparam ram_block3a12.port_a_byte_enable_clock = "none";
defparam ram_block3a12.port_a_data_out_clear = "none";
defparam ram_block3a12.port_a_data_out_clock = "none";
defparam ram_block3a12.port_a_data_width = 1;
defparam ram_block3a12.port_a_first_address = 0;
defparam ram_block3a12.port_a_first_bit_number = 12;
defparam ram_block3a12.port_a_last_address = 8191;
defparam ram_block3a12.port_a_logical_ram_depth = 16384;
defparam ram_block3a12.port_a_logical_ram_width = 32;
defparam ram_block3a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_address_clear = "none";
defparam ram_block3a12.port_b_address_clock = "clock1";
defparam ram_block3a12.port_b_address_width = 13;
defparam ram_block3a12.port_b_data_in_clock = "clock1";
defparam ram_block3a12.port_b_data_out_clear = "none";
defparam ram_block3a12.port_b_data_out_clock = "none";
defparam ram_block3a12.port_b_data_width = 1;
defparam ram_block3a12.port_b_first_address = 0;
defparam ram_block3a12.port_b_first_bit_number = 12;
defparam ram_block3a12.port_b_last_address = 8191;
defparam ram_block3a12.port_b_logical_ram_depth = 16384;
defparam ram_block3a12.port_b_logical_ram_width = 32;
defparam ram_block3a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_read_enable_clock = "clock1";
defparam ram_block3a12.port_b_write_enable_clock = "clock1";
defparam ram_block3a12.ram_block_type = "M9K";
defparam ram_block3a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014201;
// synopsys translate_on

// Location: M9K_X78_Y41_N0
cycloneive_ram_block ram_block3a45(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a45_PORTADATAOUT_bus),
	.portbdataout(ram_block3a45_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a45.clk0_core_clock_enable = "ena0";
defparam ram_block3a45.clk1_core_clock_enable = "ena1";
defparam ram_block3a45.data_interleave_offset_in_bits = 1;
defparam ram_block3a45.data_interleave_width_in_bits = 1;
defparam ram_block3a45.init_file = "meminit.hex";
defparam ram_block3a45.init_file_layout = "port_a";
defparam ram_block3a45.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a45.operation_mode = "bidir_dual_port";
defparam ram_block3a45.port_a_address_clear = "none";
defparam ram_block3a45.port_a_address_width = 13;
defparam ram_block3a45.port_a_byte_enable_clock = "none";
defparam ram_block3a45.port_a_data_out_clear = "none";
defparam ram_block3a45.port_a_data_out_clock = "none";
defparam ram_block3a45.port_a_data_width = 1;
defparam ram_block3a45.port_a_first_address = 0;
defparam ram_block3a45.port_a_first_bit_number = 13;
defparam ram_block3a45.port_a_last_address = 8191;
defparam ram_block3a45.port_a_logical_ram_depth = 16384;
defparam ram_block3a45.port_a_logical_ram_width = 32;
defparam ram_block3a45.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_address_clear = "none";
defparam ram_block3a45.port_b_address_clock = "clock1";
defparam ram_block3a45.port_b_address_width = 13;
defparam ram_block3a45.port_b_data_in_clock = "clock1";
defparam ram_block3a45.port_b_data_out_clear = "none";
defparam ram_block3a45.port_b_data_out_clock = "none";
defparam ram_block3a45.port_b_data_width = 1;
defparam ram_block3a45.port_b_first_address = 0;
defparam ram_block3a45.port_b_first_bit_number = 13;
defparam ram_block3a45.port_b_last_address = 8191;
defparam ram_block3a45.port_b_logical_ram_depth = 16384;
defparam ram_block3a45.port_b_logical_ram_width = 32;
defparam ram_block3a45.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_read_enable_clock = "clock1";
defparam ram_block3a45.port_b_write_enable_clock = "clock1";
defparam ram_block3a45.ram_block_type = "M9K";
defparam ram_block3a45.mem_init3 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001F9FD388D4AF84D1421FCDE7200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y43_N0
cycloneive_ram_block ram_block3a13(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a13_PORTADATAOUT_bus),
	.portbdataout(ram_block3a13_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a13.clk0_core_clock_enable = "ena0";
defparam ram_block3a13.clk1_core_clock_enable = "ena1";
defparam ram_block3a13.data_interleave_offset_in_bits = 1;
defparam ram_block3a13.data_interleave_width_in_bits = 1;
defparam ram_block3a13.init_file = "meminit.hex";
defparam ram_block3a13.init_file_layout = "port_a";
defparam ram_block3a13.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a13.operation_mode = "bidir_dual_port";
defparam ram_block3a13.port_a_address_clear = "none";
defparam ram_block3a13.port_a_address_width = 13;
defparam ram_block3a13.port_a_byte_enable_clock = "none";
defparam ram_block3a13.port_a_data_out_clear = "none";
defparam ram_block3a13.port_a_data_out_clock = "none";
defparam ram_block3a13.port_a_data_width = 1;
defparam ram_block3a13.port_a_first_address = 0;
defparam ram_block3a13.port_a_first_bit_number = 13;
defparam ram_block3a13.port_a_last_address = 8191;
defparam ram_block3a13.port_a_logical_ram_depth = 16384;
defparam ram_block3a13.port_a_logical_ram_width = 32;
defparam ram_block3a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_address_clear = "none";
defparam ram_block3a13.port_b_address_clock = "clock1";
defparam ram_block3a13.port_b_address_width = 13;
defparam ram_block3a13.port_b_data_in_clock = "clock1";
defparam ram_block3a13.port_b_data_out_clear = "none";
defparam ram_block3a13.port_b_data_out_clock = "none";
defparam ram_block3a13.port_b_data_width = 1;
defparam ram_block3a13.port_b_first_address = 0;
defparam ram_block3a13.port_b_first_bit_number = 13;
defparam ram_block3a13.port_b_last_address = 8191;
defparam ram_block3a13.port_b_logical_ram_depth = 16384;
defparam ram_block3a13.port_b_logical_ram_width = 32;
defparam ram_block3a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_read_enable_clock = "clock1";
defparam ram_block3a13.port_b_write_enable_clock = "clock1";
defparam ram_block3a13.ram_block_type = "M9K";
defparam ram_block3a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000015A01;
// synopsys translate_on

// Location: M9K_X78_Y32_N0
cycloneive_ram_block ram_block3a46(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a46_PORTADATAOUT_bus),
	.portbdataout(ram_block3a46_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a46.clk0_core_clock_enable = "ena0";
defparam ram_block3a46.clk1_core_clock_enable = "ena1";
defparam ram_block3a46.data_interleave_offset_in_bits = 1;
defparam ram_block3a46.data_interleave_width_in_bits = 1;
defparam ram_block3a46.init_file = "meminit.hex";
defparam ram_block3a46.init_file_layout = "port_a";
defparam ram_block3a46.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a46.operation_mode = "bidir_dual_port";
defparam ram_block3a46.port_a_address_clear = "none";
defparam ram_block3a46.port_a_address_width = 13;
defparam ram_block3a46.port_a_byte_enable_clock = "none";
defparam ram_block3a46.port_a_data_out_clear = "none";
defparam ram_block3a46.port_a_data_out_clock = "none";
defparam ram_block3a46.port_a_data_width = 1;
defparam ram_block3a46.port_a_first_address = 0;
defparam ram_block3a46.port_a_first_bit_number = 14;
defparam ram_block3a46.port_a_last_address = 8191;
defparam ram_block3a46.port_a_logical_ram_depth = 16384;
defparam ram_block3a46.port_a_logical_ram_width = 32;
defparam ram_block3a46.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_address_clear = "none";
defparam ram_block3a46.port_b_address_clock = "clock1";
defparam ram_block3a46.port_b_address_width = 13;
defparam ram_block3a46.port_b_data_in_clock = "clock1";
defparam ram_block3a46.port_b_data_out_clear = "none";
defparam ram_block3a46.port_b_data_out_clock = "none";
defparam ram_block3a46.port_b_data_width = 1;
defparam ram_block3a46.port_b_first_address = 0;
defparam ram_block3a46.port_b_first_bit_number = 14;
defparam ram_block3a46.port_b_last_address = 8191;
defparam ram_block3a46.port_b_logical_ram_depth = 16384;
defparam ram_block3a46.port_b_logical_ram_width = 32;
defparam ram_block3a46.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_read_enable_clock = "clock1";
defparam ram_block3a46.port_b_write_enable_clock = "clock1";
defparam ram_block3a46.ram_block_type = "M9K";
defparam ram_block3a46.mem_init3 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006016FF21E8A5086CEC071A7D20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y33_N0
cycloneive_ram_block ram_block3a14(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a14_PORTADATAOUT_bus),
	.portbdataout(ram_block3a14_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a14.clk0_core_clock_enable = "ena0";
defparam ram_block3a14.clk1_core_clock_enable = "ena1";
defparam ram_block3a14.data_interleave_offset_in_bits = 1;
defparam ram_block3a14.data_interleave_width_in_bits = 1;
defparam ram_block3a14.init_file = "meminit.hex";
defparam ram_block3a14.init_file_layout = "port_a";
defparam ram_block3a14.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a14.operation_mode = "bidir_dual_port";
defparam ram_block3a14.port_a_address_clear = "none";
defparam ram_block3a14.port_a_address_width = 13;
defparam ram_block3a14.port_a_byte_enable_clock = "none";
defparam ram_block3a14.port_a_data_out_clear = "none";
defparam ram_block3a14.port_a_data_out_clock = "none";
defparam ram_block3a14.port_a_data_width = 1;
defparam ram_block3a14.port_a_first_address = 0;
defparam ram_block3a14.port_a_first_bit_number = 14;
defparam ram_block3a14.port_a_last_address = 8191;
defparam ram_block3a14.port_a_logical_ram_depth = 16384;
defparam ram_block3a14.port_a_logical_ram_width = 32;
defparam ram_block3a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_address_clear = "none";
defparam ram_block3a14.port_b_address_clock = "clock1";
defparam ram_block3a14.port_b_address_width = 13;
defparam ram_block3a14.port_b_data_in_clock = "clock1";
defparam ram_block3a14.port_b_data_out_clear = "none";
defparam ram_block3a14.port_b_data_out_clock = "none";
defparam ram_block3a14.port_b_data_width = 1;
defparam ram_block3a14.port_b_first_address = 0;
defparam ram_block3a14.port_b_first_bit_number = 14;
defparam ram_block3a14.port_b_last_address = 8191;
defparam ram_block3a14.port_b_logical_ram_depth = 16384;
defparam ram_block3a14.port_b_logical_ram_width = 32;
defparam ram_block3a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_read_enable_clock = "clock1";
defparam ram_block3a14.port_b_write_enable_clock = "clock1";
defparam ram_block3a14.ram_block_type = "M9K";
defparam ram_block3a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014001;
// synopsys translate_on

// Location: M9K_X78_Y42_N0
cycloneive_ram_block ram_block3a47(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a47_PORTADATAOUT_bus),
	.portbdataout(ram_block3a47_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a47.clk0_core_clock_enable = "ena0";
defparam ram_block3a47.clk1_core_clock_enable = "ena1";
defparam ram_block3a47.data_interleave_offset_in_bits = 1;
defparam ram_block3a47.data_interleave_width_in_bits = 1;
defparam ram_block3a47.init_file = "meminit.hex";
defparam ram_block3a47.init_file_layout = "port_a";
defparam ram_block3a47.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a47.operation_mode = "bidir_dual_port";
defparam ram_block3a47.port_a_address_clear = "none";
defparam ram_block3a47.port_a_address_width = 13;
defparam ram_block3a47.port_a_byte_enable_clock = "none";
defparam ram_block3a47.port_a_data_out_clear = "none";
defparam ram_block3a47.port_a_data_out_clock = "none";
defparam ram_block3a47.port_a_data_width = 1;
defparam ram_block3a47.port_a_first_address = 0;
defparam ram_block3a47.port_a_first_bit_number = 15;
defparam ram_block3a47.port_a_last_address = 8191;
defparam ram_block3a47.port_a_logical_ram_depth = 16384;
defparam ram_block3a47.port_a_logical_ram_width = 32;
defparam ram_block3a47.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_address_clear = "none";
defparam ram_block3a47.port_b_address_clock = "clock1";
defparam ram_block3a47.port_b_address_width = 13;
defparam ram_block3a47.port_b_data_in_clock = "clock1";
defparam ram_block3a47.port_b_data_out_clear = "none";
defparam ram_block3a47.port_b_data_out_clock = "none";
defparam ram_block3a47.port_b_data_width = 1;
defparam ram_block3a47.port_b_first_address = 0;
defparam ram_block3a47.port_b_first_bit_number = 15;
defparam ram_block3a47.port_b_last_address = 8191;
defparam ram_block3a47.port_b_logical_ram_depth = 16384;
defparam ram_block3a47.port_b_logical_ram_width = 32;
defparam ram_block3a47.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_read_enable_clock = "clock1";
defparam ram_block3a47.port_b_write_enable_clock = "clock1";
defparam ram_block3a47.ram_block_type = "M9K";
defparam ram_block3a47.mem_init3 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FEF9FF77AC95FDC4AE96A58200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y42_N0
cycloneive_ram_block ram_block3a15(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a15_PORTADATAOUT_bus),
	.portbdataout(ram_block3a15_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a15.clk0_core_clock_enable = "ena0";
defparam ram_block3a15.clk1_core_clock_enable = "ena1";
defparam ram_block3a15.data_interleave_offset_in_bits = 1;
defparam ram_block3a15.data_interleave_width_in_bits = 1;
defparam ram_block3a15.init_file = "meminit.hex";
defparam ram_block3a15.init_file_layout = "port_a";
defparam ram_block3a15.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a15.operation_mode = "bidir_dual_port";
defparam ram_block3a15.port_a_address_clear = "none";
defparam ram_block3a15.port_a_address_width = 13;
defparam ram_block3a15.port_a_byte_enable_clock = "none";
defparam ram_block3a15.port_a_data_out_clear = "none";
defparam ram_block3a15.port_a_data_out_clock = "none";
defparam ram_block3a15.port_a_data_width = 1;
defparam ram_block3a15.port_a_first_address = 0;
defparam ram_block3a15.port_a_first_bit_number = 15;
defparam ram_block3a15.port_a_last_address = 8191;
defparam ram_block3a15.port_a_logical_ram_depth = 16384;
defparam ram_block3a15.port_a_logical_ram_width = 32;
defparam ram_block3a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_address_clear = "none";
defparam ram_block3a15.port_b_address_clock = "clock1";
defparam ram_block3a15.port_b_address_width = 13;
defparam ram_block3a15.port_b_data_in_clock = "clock1";
defparam ram_block3a15.port_b_data_out_clear = "none";
defparam ram_block3a15.port_b_data_out_clock = "none";
defparam ram_block3a15.port_b_data_width = 1;
defparam ram_block3a15.port_b_first_address = 0;
defparam ram_block3a15.port_b_first_bit_number = 15;
defparam ram_block3a15.port_b_last_address = 8191;
defparam ram_block3a15.port_b_logical_ram_depth = 16384;
defparam ram_block3a15.port_b_logical_ram_width = 32;
defparam ram_block3a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_read_enable_clock = "clock1";
defparam ram_block3a15.port_b_write_enable_clock = "clock1";
defparam ram_block3a15.ram_block_type = "M9K";
defparam ram_block3a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014001;
// synopsys translate_on

// Location: M9K_X78_Y44_N0
cycloneive_ram_block ram_block3a48(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a48_PORTADATAOUT_bus),
	.portbdataout(ram_block3a48_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a48.clk0_core_clock_enable = "ena0";
defparam ram_block3a48.clk1_core_clock_enable = "ena1";
defparam ram_block3a48.data_interleave_offset_in_bits = 1;
defparam ram_block3a48.data_interleave_width_in_bits = 1;
defparam ram_block3a48.init_file = "meminit.hex";
defparam ram_block3a48.init_file_layout = "port_a";
defparam ram_block3a48.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a48.operation_mode = "bidir_dual_port";
defparam ram_block3a48.port_a_address_clear = "none";
defparam ram_block3a48.port_a_address_width = 13;
defparam ram_block3a48.port_a_byte_enable_clock = "none";
defparam ram_block3a48.port_a_data_out_clear = "none";
defparam ram_block3a48.port_a_data_out_clock = "none";
defparam ram_block3a48.port_a_data_width = 1;
defparam ram_block3a48.port_a_first_address = 0;
defparam ram_block3a48.port_a_first_bit_number = 16;
defparam ram_block3a48.port_a_last_address = 8191;
defparam ram_block3a48.port_a_logical_ram_depth = 16384;
defparam ram_block3a48.port_a_logical_ram_width = 32;
defparam ram_block3a48.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_address_clear = "none";
defparam ram_block3a48.port_b_address_clock = "clock1";
defparam ram_block3a48.port_b_address_width = 13;
defparam ram_block3a48.port_b_data_in_clock = "clock1";
defparam ram_block3a48.port_b_data_out_clear = "none";
defparam ram_block3a48.port_b_data_out_clock = "none";
defparam ram_block3a48.port_b_data_width = 1;
defparam ram_block3a48.port_b_first_address = 0;
defparam ram_block3a48.port_b_first_bit_number = 16;
defparam ram_block3a48.port_b_last_address = 8191;
defparam ram_block3a48.port_b_logical_ram_depth = 16384;
defparam ram_block3a48.port_b_logical_ram_width = 32;
defparam ram_block3a48.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_read_enable_clock = "clock1";
defparam ram_block3a48.port_b_write_enable_clock = "clock1";
defparam ram_block3a48.ram_block_type = "M9K";
defparam ram_block3a48.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y46_N0
cycloneive_ram_block ram_block3a16(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a16_PORTADATAOUT_bus),
	.portbdataout(ram_block3a16_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a16.clk0_core_clock_enable = "ena0";
defparam ram_block3a16.clk1_core_clock_enable = "ena1";
defparam ram_block3a16.data_interleave_offset_in_bits = 1;
defparam ram_block3a16.data_interleave_width_in_bits = 1;
defparam ram_block3a16.init_file = "meminit.hex";
defparam ram_block3a16.init_file_layout = "port_a";
defparam ram_block3a16.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a16.operation_mode = "bidir_dual_port";
defparam ram_block3a16.port_a_address_clear = "none";
defparam ram_block3a16.port_a_address_width = 13;
defparam ram_block3a16.port_a_byte_enable_clock = "none";
defparam ram_block3a16.port_a_data_out_clear = "none";
defparam ram_block3a16.port_a_data_out_clock = "none";
defparam ram_block3a16.port_a_data_width = 1;
defparam ram_block3a16.port_a_first_address = 0;
defparam ram_block3a16.port_a_first_bit_number = 16;
defparam ram_block3a16.port_a_last_address = 8191;
defparam ram_block3a16.port_a_logical_ram_depth = 16384;
defparam ram_block3a16.port_a_logical_ram_width = 32;
defparam ram_block3a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_address_clear = "none";
defparam ram_block3a16.port_b_address_clock = "clock1";
defparam ram_block3a16.port_b_address_width = 13;
defparam ram_block3a16.port_b_data_in_clock = "clock1";
defparam ram_block3a16.port_b_data_out_clear = "none";
defparam ram_block3a16.port_b_data_out_clock = "none";
defparam ram_block3a16.port_b_data_width = 1;
defparam ram_block3a16.port_b_first_address = 0;
defparam ram_block3a16.port_b_first_bit_number = 16;
defparam ram_block3a16.port_b_last_address = 8191;
defparam ram_block3a16.port_b_logical_ram_depth = 16384;
defparam ram_block3a16.port_b_logical_ram_width = 32;
defparam ram_block3a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_read_enable_clock = "clock1";
defparam ram_block3a16.port_b_write_enable_clock = "clock1";
defparam ram_block3a16.ram_block_type = "M9K";
defparam ram_block3a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000019253;
// synopsys translate_on

// Location: M9K_X37_Y43_N0
cycloneive_ram_block ram_block3a49(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a49_PORTADATAOUT_bus),
	.portbdataout(ram_block3a49_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a49.clk0_core_clock_enable = "ena0";
defparam ram_block3a49.clk1_core_clock_enable = "ena1";
defparam ram_block3a49.data_interleave_offset_in_bits = 1;
defparam ram_block3a49.data_interleave_width_in_bits = 1;
defparam ram_block3a49.init_file = "meminit.hex";
defparam ram_block3a49.init_file_layout = "port_a";
defparam ram_block3a49.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a49.operation_mode = "bidir_dual_port";
defparam ram_block3a49.port_a_address_clear = "none";
defparam ram_block3a49.port_a_address_width = 13;
defparam ram_block3a49.port_a_byte_enable_clock = "none";
defparam ram_block3a49.port_a_data_out_clear = "none";
defparam ram_block3a49.port_a_data_out_clock = "none";
defparam ram_block3a49.port_a_data_width = 1;
defparam ram_block3a49.port_a_first_address = 0;
defparam ram_block3a49.port_a_first_bit_number = 17;
defparam ram_block3a49.port_a_last_address = 8191;
defparam ram_block3a49.port_a_logical_ram_depth = 16384;
defparam ram_block3a49.port_a_logical_ram_width = 32;
defparam ram_block3a49.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_address_clear = "none";
defparam ram_block3a49.port_b_address_clock = "clock1";
defparam ram_block3a49.port_b_address_width = 13;
defparam ram_block3a49.port_b_data_in_clock = "clock1";
defparam ram_block3a49.port_b_data_out_clear = "none";
defparam ram_block3a49.port_b_data_out_clock = "none";
defparam ram_block3a49.port_b_data_width = 1;
defparam ram_block3a49.port_b_first_address = 0;
defparam ram_block3a49.port_b_first_bit_number = 17;
defparam ram_block3a49.port_b_last_address = 8191;
defparam ram_block3a49.port_b_logical_ram_depth = 16384;
defparam ram_block3a49.port_b_logical_ram_width = 32;
defparam ram_block3a49.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_read_enable_clock = "clock1";
defparam ram_block3a49.port_b_write_enable_clock = "clock1";
defparam ram_block3a49.ram_block_type = "M9K";
defparam ram_block3a49.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y44_N0
cycloneive_ram_block ram_block3a17(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a17_PORTADATAOUT_bus),
	.portbdataout(ram_block3a17_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a17.clk0_core_clock_enable = "ena0";
defparam ram_block3a17.clk1_core_clock_enable = "ena1";
defparam ram_block3a17.data_interleave_offset_in_bits = 1;
defparam ram_block3a17.data_interleave_width_in_bits = 1;
defparam ram_block3a17.init_file = "meminit.hex";
defparam ram_block3a17.init_file_layout = "port_a";
defparam ram_block3a17.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a17.operation_mode = "bidir_dual_port";
defparam ram_block3a17.port_a_address_clear = "none";
defparam ram_block3a17.port_a_address_width = 13;
defparam ram_block3a17.port_a_byte_enable_clock = "none";
defparam ram_block3a17.port_a_data_out_clear = "none";
defparam ram_block3a17.port_a_data_out_clock = "none";
defparam ram_block3a17.port_a_data_width = 1;
defparam ram_block3a17.port_a_first_address = 0;
defparam ram_block3a17.port_a_first_bit_number = 17;
defparam ram_block3a17.port_a_last_address = 8191;
defparam ram_block3a17.port_a_logical_ram_depth = 16384;
defparam ram_block3a17.port_a_logical_ram_width = 32;
defparam ram_block3a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_address_clear = "none";
defparam ram_block3a17.port_b_address_clock = "clock1";
defparam ram_block3a17.port_b_address_width = 13;
defparam ram_block3a17.port_b_data_in_clock = "clock1";
defparam ram_block3a17.port_b_data_out_clear = "none";
defparam ram_block3a17.port_b_data_out_clock = "none";
defparam ram_block3a17.port_b_data_width = 1;
defparam ram_block3a17.port_b_first_address = 0;
defparam ram_block3a17.port_b_first_bit_number = 17;
defparam ram_block3a17.port_b_last_address = 8191;
defparam ram_block3a17.port_b_logical_ram_depth = 16384;
defparam ram_block3a17.port_b_logical_ram_width = 32;
defparam ram_block3a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_read_enable_clock = "clock1";
defparam ram_block3a17.port_b_write_enable_clock = "clock1";
defparam ram_block3a17.ram_block_type = "M9K";
defparam ram_block3a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010A94;
// synopsys translate_on

// Location: M9K_X64_Y45_N0
cycloneive_ram_block ram_block3a50(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a50_PORTADATAOUT_bus),
	.portbdataout(ram_block3a50_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a50.clk0_core_clock_enable = "ena0";
defparam ram_block3a50.clk1_core_clock_enable = "ena1";
defparam ram_block3a50.data_interleave_offset_in_bits = 1;
defparam ram_block3a50.data_interleave_width_in_bits = 1;
defparam ram_block3a50.init_file = "meminit.hex";
defparam ram_block3a50.init_file_layout = "port_a";
defparam ram_block3a50.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a50.operation_mode = "bidir_dual_port";
defparam ram_block3a50.port_a_address_clear = "none";
defparam ram_block3a50.port_a_address_width = 13;
defparam ram_block3a50.port_a_byte_enable_clock = "none";
defparam ram_block3a50.port_a_data_out_clear = "none";
defparam ram_block3a50.port_a_data_out_clock = "none";
defparam ram_block3a50.port_a_data_width = 1;
defparam ram_block3a50.port_a_first_address = 0;
defparam ram_block3a50.port_a_first_bit_number = 18;
defparam ram_block3a50.port_a_last_address = 8191;
defparam ram_block3a50.port_a_logical_ram_depth = 16384;
defparam ram_block3a50.port_a_logical_ram_width = 32;
defparam ram_block3a50.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_address_clear = "none";
defparam ram_block3a50.port_b_address_clock = "clock1";
defparam ram_block3a50.port_b_address_width = 13;
defparam ram_block3a50.port_b_data_in_clock = "clock1";
defparam ram_block3a50.port_b_data_out_clear = "none";
defparam ram_block3a50.port_b_data_out_clock = "none";
defparam ram_block3a50.port_b_data_width = 1;
defparam ram_block3a50.port_b_first_address = 0;
defparam ram_block3a50.port_b_first_bit_number = 18;
defparam ram_block3a50.port_b_last_address = 8191;
defparam ram_block3a50.port_b_logical_ram_depth = 16384;
defparam ram_block3a50.port_b_logical_ram_width = 32;
defparam ram_block3a50.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_read_enable_clock = "clock1";
defparam ram_block3a50.port_b_write_enable_clock = "clock1";
defparam ram_block3a50.ram_block_type = "M9K";
defparam ram_block3a50.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y46_N0
cycloneive_ram_block ram_block3a18(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a18_PORTADATAOUT_bus),
	.portbdataout(ram_block3a18_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a18.clk0_core_clock_enable = "ena0";
defparam ram_block3a18.clk1_core_clock_enable = "ena1";
defparam ram_block3a18.data_interleave_offset_in_bits = 1;
defparam ram_block3a18.data_interleave_width_in_bits = 1;
defparam ram_block3a18.init_file = "meminit.hex";
defparam ram_block3a18.init_file_layout = "port_a";
defparam ram_block3a18.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a18.operation_mode = "bidir_dual_port";
defparam ram_block3a18.port_a_address_clear = "none";
defparam ram_block3a18.port_a_address_width = 13;
defparam ram_block3a18.port_a_byte_enable_clock = "none";
defparam ram_block3a18.port_a_data_out_clear = "none";
defparam ram_block3a18.port_a_data_out_clock = "none";
defparam ram_block3a18.port_a_data_width = 1;
defparam ram_block3a18.port_a_first_address = 0;
defparam ram_block3a18.port_a_first_bit_number = 18;
defparam ram_block3a18.port_a_last_address = 8191;
defparam ram_block3a18.port_a_logical_ram_depth = 16384;
defparam ram_block3a18.port_a_logical_ram_width = 32;
defparam ram_block3a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_address_clear = "none";
defparam ram_block3a18.port_b_address_clock = "clock1";
defparam ram_block3a18.port_b_address_width = 13;
defparam ram_block3a18.port_b_data_in_clock = "clock1";
defparam ram_block3a18.port_b_data_out_clear = "none";
defparam ram_block3a18.port_b_data_out_clock = "none";
defparam ram_block3a18.port_b_data_width = 1;
defparam ram_block3a18.port_b_first_address = 0;
defparam ram_block3a18.port_b_first_bit_number = 18;
defparam ram_block3a18.port_b_last_address = 8191;
defparam ram_block3a18.port_b_logical_ram_depth = 16384;
defparam ram_block3a18.port_b_logical_ram_width = 32;
defparam ram_block3a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_read_enable_clock = "clock1";
defparam ram_block3a18.port_b_write_enable_clock = "clock1";
defparam ram_block3a18.ram_block_type = "M9K";
defparam ram_block3a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000180E1;
// synopsys translate_on

// Location: M9K_X51_Y43_N0
cycloneive_ram_block ram_block3a51(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a51_PORTADATAOUT_bus),
	.portbdataout(ram_block3a51_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a51.clk0_core_clock_enable = "ena0";
defparam ram_block3a51.clk1_core_clock_enable = "ena1";
defparam ram_block3a51.data_interleave_offset_in_bits = 1;
defparam ram_block3a51.data_interleave_width_in_bits = 1;
defparam ram_block3a51.init_file = "meminit.hex";
defparam ram_block3a51.init_file_layout = "port_a";
defparam ram_block3a51.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a51.operation_mode = "bidir_dual_port";
defparam ram_block3a51.port_a_address_clear = "none";
defparam ram_block3a51.port_a_address_width = 13;
defparam ram_block3a51.port_a_byte_enable_clock = "none";
defparam ram_block3a51.port_a_data_out_clear = "none";
defparam ram_block3a51.port_a_data_out_clock = "none";
defparam ram_block3a51.port_a_data_width = 1;
defparam ram_block3a51.port_a_first_address = 0;
defparam ram_block3a51.port_a_first_bit_number = 19;
defparam ram_block3a51.port_a_last_address = 8191;
defparam ram_block3a51.port_a_logical_ram_depth = 16384;
defparam ram_block3a51.port_a_logical_ram_width = 32;
defparam ram_block3a51.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_address_clear = "none";
defparam ram_block3a51.port_b_address_clock = "clock1";
defparam ram_block3a51.port_b_address_width = 13;
defparam ram_block3a51.port_b_data_in_clock = "clock1";
defparam ram_block3a51.port_b_data_out_clear = "none";
defparam ram_block3a51.port_b_data_out_clock = "none";
defparam ram_block3a51.port_b_data_width = 1;
defparam ram_block3a51.port_b_first_address = 0;
defparam ram_block3a51.port_b_first_bit_number = 19;
defparam ram_block3a51.port_b_last_address = 8191;
defparam ram_block3a51.port_b_logical_ram_depth = 16384;
defparam ram_block3a51.port_b_logical_ram_width = 32;
defparam ram_block3a51.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_read_enable_clock = "clock1";
defparam ram_block3a51.port_b_write_enable_clock = "clock1";
defparam ram_block3a51.ram_block_type = "M9K";
defparam ram_block3a51.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y38_N0
cycloneive_ram_block ram_block3a19(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a19_PORTADATAOUT_bus),
	.portbdataout(ram_block3a19_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a19.clk0_core_clock_enable = "ena0";
defparam ram_block3a19.clk1_core_clock_enable = "ena1";
defparam ram_block3a19.data_interleave_offset_in_bits = 1;
defparam ram_block3a19.data_interleave_width_in_bits = 1;
defparam ram_block3a19.init_file = "meminit.hex";
defparam ram_block3a19.init_file_layout = "port_a";
defparam ram_block3a19.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a19.operation_mode = "bidir_dual_port";
defparam ram_block3a19.port_a_address_clear = "none";
defparam ram_block3a19.port_a_address_width = 13;
defparam ram_block3a19.port_a_byte_enable_clock = "none";
defparam ram_block3a19.port_a_data_out_clear = "none";
defparam ram_block3a19.port_a_data_out_clock = "none";
defparam ram_block3a19.port_a_data_width = 1;
defparam ram_block3a19.port_a_first_address = 0;
defparam ram_block3a19.port_a_first_bit_number = 19;
defparam ram_block3a19.port_a_last_address = 8191;
defparam ram_block3a19.port_a_logical_ram_depth = 16384;
defparam ram_block3a19.port_a_logical_ram_width = 32;
defparam ram_block3a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_address_clear = "none";
defparam ram_block3a19.port_b_address_clock = "clock1";
defparam ram_block3a19.port_b_address_width = 13;
defparam ram_block3a19.port_b_data_in_clock = "clock1";
defparam ram_block3a19.port_b_data_out_clear = "none";
defparam ram_block3a19.port_b_data_out_clock = "none";
defparam ram_block3a19.port_b_data_width = 1;
defparam ram_block3a19.port_b_first_address = 0;
defparam ram_block3a19.port_b_first_bit_number = 19;
defparam ram_block3a19.port_b_last_address = 8191;
defparam ram_block3a19.port_b_logical_ram_depth = 16384;
defparam ram_block3a19.port_b_logical_ram_width = 32;
defparam ram_block3a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_read_enable_clock = "clock1";
defparam ram_block3a19.port_b_write_enable_clock = "clock1";
defparam ram_block3a19.ram_block_type = "M9K";
defparam ram_block3a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001;
// synopsys translate_on

// Location: M9K_X64_Y31_N0
cycloneive_ram_block ram_block3a52(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a52_PORTADATAOUT_bus),
	.portbdataout(ram_block3a52_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a52.clk0_core_clock_enable = "ena0";
defparam ram_block3a52.clk1_core_clock_enable = "ena1";
defparam ram_block3a52.data_interleave_offset_in_bits = 1;
defparam ram_block3a52.data_interleave_width_in_bits = 1;
defparam ram_block3a52.init_file = "meminit.hex";
defparam ram_block3a52.init_file_layout = "port_a";
defparam ram_block3a52.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a52.operation_mode = "bidir_dual_port";
defparam ram_block3a52.port_a_address_clear = "none";
defparam ram_block3a52.port_a_address_width = 13;
defparam ram_block3a52.port_a_byte_enable_clock = "none";
defparam ram_block3a52.port_a_data_out_clear = "none";
defparam ram_block3a52.port_a_data_out_clock = "none";
defparam ram_block3a52.port_a_data_width = 1;
defparam ram_block3a52.port_a_first_address = 0;
defparam ram_block3a52.port_a_first_bit_number = 20;
defparam ram_block3a52.port_a_last_address = 8191;
defparam ram_block3a52.port_a_logical_ram_depth = 16384;
defparam ram_block3a52.port_a_logical_ram_width = 32;
defparam ram_block3a52.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_address_clear = "none";
defparam ram_block3a52.port_b_address_clock = "clock1";
defparam ram_block3a52.port_b_address_width = 13;
defparam ram_block3a52.port_b_data_in_clock = "clock1";
defparam ram_block3a52.port_b_data_out_clear = "none";
defparam ram_block3a52.port_b_data_out_clock = "none";
defparam ram_block3a52.port_b_data_width = 1;
defparam ram_block3a52.port_b_first_address = 0;
defparam ram_block3a52.port_b_first_bit_number = 20;
defparam ram_block3a52.port_b_last_address = 8191;
defparam ram_block3a52.port_b_logical_ram_depth = 16384;
defparam ram_block3a52.port_b_logical_ram_width = 32;
defparam ram_block3a52.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_read_enable_clock = "clock1";
defparam ram_block3a52.port_b_write_enable_clock = "clock1";
defparam ram_block3a52.ram_block_type = "M9K";
defparam ram_block3a52.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y35_N0
cycloneive_ram_block ram_block3a20(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a20_PORTADATAOUT_bus),
	.portbdataout(ram_block3a20_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a20.clk0_core_clock_enable = "ena0";
defparam ram_block3a20.clk1_core_clock_enable = "ena1";
defparam ram_block3a20.data_interleave_offset_in_bits = 1;
defparam ram_block3a20.data_interleave_width_in_bits = 1;
defparam ram_block3a20.init_file = "meminit.hex";
defparam ram_block3a20.init_file_layout = "port_a";
defparam ram_block3a20.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a20.operation_mode = "bidir_dual_port";
defparam ram_block3a20.port_a_address_clear = "none";
defparam ram_block3a20.port_a_address_width = 13;
defparam ram_block3a20.port_a_byte_enable_clock = "none";
defparam ram_block3a20.port_a_data_out_clear = "none";
defparam ram_block3a20.port_a_data_out_clock = "none";
defparam ram_block3a20.port_a_data_width = 1;
defparam ram_block3a20.port_a_first_address = 0;
defparam ram_block3a20.port_a_first_bit_number = 20;
defparam ram_block3a20.port_a_last_address = 8191;
defparam ram_block3a20.port_a_logical_ram_depth = 16384;
defparam ram_block3a20.port_a_logical_ram_width = 32;
defparam ram_block3a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_address_clear = "none";
defparam ram_block3a20.port_b_address_clock = "clock1";
defparam ram_block3a20.port_b_address_width = 13;
defparam ram_block3a20.port_b_data_in_clock = "clock1";
defparam ram_block3a20.port_b_data_out_clear = "none";
defparam ram_block3a20.port_b_data_out_clock = "none";
defparam ram_block3a20.port_b_data_width = 1;
defparam ram_block3a20.port_b_first_address = 0;
defparam ram_block3a20.port_b_first_bit_number = 20;
defparam ram_block3a20.port_b_last_address = 8191;
defparam ram_block3a20.port_b_logical_ram_depth = 16384;
defparam ram_block3a20.port_b_logical_ram_width = 32;
defparam ram_block3a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_read_enable_clock = "clock1";
defparam ram_block3a20.port_b_write_enable_clock = "clock1";
defparam ram_block3a20.ram_block_type = "M9K";
defparam ram_block3a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001;
// synopsys translate_on

// Location: M9K_X37_Y37_N0
cycloneive_ram_block ram_block3a53(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a53_PORTADATAOUT_bus),
	.portbdataout(ram_block3a53_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a53.clk0_core_clock_enable = "ena0";
defparam ram_block3a53.clk1_core_clock_enable = "ena1";
defparam ram_block3a53.data_interleave_offset_in_bits = 1;
defparam ram_block3a53.data_interleave_width_in_bits = 1;
defparam ram_block3a53.init_file = "meminit.hex";
defparam ram_block3a53.init_file_layout = "port_a";
defparam ram_block3a53.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a53.operation_mode = "bidir_dual_port";
defparam ram_block3a53.port_a_address_clear = "none";
defparam ram_block3a53.port_a_address_width = 13;
defparam ram_block3a53.port_a_byte_enable_clock = "none";
defparam ram_block3a53.port_a_data_out_clear = "none";
defparam ram_block3a53.port_a_data_out_clock = "none";
defparam ram_block3a53.port_a_data_width = 1;
defparam ram_block3a53.port_a_first_address = 0;
defparam ram_block3a53.port_a_first_bit_number = 21;
defparam ram_block3a53.port_a_last_address = 8191;
defparam ram_block3a53.port_a_logical_ram_depth = 16384;
defparam ram_block3a53.port_a_logical_ram_width = 32;
defparam ram_block3a53.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_address_clear = "none";
defparam ram_block3a53.port_b_address_clock = "clock1";
defparam ram_block3a53.port_b_address_width = 13;
defparam ram_block3a53.port_b_data_in_clock = "clock1";
defparam ram_block3a53.port_b_data_out_clear = "none";
defparam ram_block3a53.port_b_data_out_clock = "none";
defparam ram_block3a53.port_b_data_width = 1;
defparam ram_block3a53.port_b_first_address = 0;
defparam ram_block3a53.port_b_first_bit_number = 21;
defparam ram_block3a53.port_b_last_address = 8191;
defparam ram_block3a53.port_b_logical_ram_depth = 16384;
defparam ram_block3a53.port_b_logical_ram_width = 32;
defparam ram_block3a53.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_read_enable_clock = "clock1";
defparam ram_block3a53.port_b_write_enable_clock = "clock1";
defparam ram_block3a53.ram_block_type = "M9K";
defparam ram_block3a53.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y39_N0
cycloneive_ram_block ram_block3a21(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a21_PORTADATAOUT_bus),
	.portbdataout(ram_block3a21_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a21.clk0_core_clock_enable = "ena0";
defparam ram_block3a21.clk1_core_clock_enable = "ena1";
defparam ram_block3a21.data_interleave_offset_in_bits = 1;
defparam ram_block3a21.data_interleave_width_in_bits = 1;
defparam ram_block3a21.init_file = "meminit.hex";
defparam ram_block3a21.init_file_layout = "port_a";
defparam ram_block3a21.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a21.operation_mode = "bidir_dual_port";
defparam ram_block3a21.port_a_address_clear = "none";
defparam ram_block3a21.port_a_address_width = 13;
defparam ram_block3a21.port_a_byte_enable_clock = "none";
defparam ram_block3a21.port_a_data_out_clear = "none";
defparam ram_block3a21.port_a_data_out_clock = "none";
defparam ram_block3a21.port_a_data_width = 1;
defparam ram_block3a21.port_a_first_address = 0;
defparam ram_block3a21.port_a_first_bit_number = 21;
defparam ram_block3a21.port_a_last_address = 8191;
defparam ram_block3a21.port_a_logical_ram_depth = 16384;
defparam ram_block3a21.port_a_logical_ram_width = 32;
defparam ram_block3a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_address_clear = "none";
defparam ram_block3a21.port_b_address_clock = "clock1";
defparam ram_block3a21.port_b_address_width = 13;
defparam ram_block3a21.port_b_data_in_clock = "clock1";
defparam ram_block3a21.port_b_data_out_clear = "none";
defparam ram_block3a21.port_b_data_out_clock = "none";
defparam ram_block3a21.port_b_data_width = 1;
defparam ram_block3a21.port_b_first_address = 0;
defparam ram_block3a21.port_b_first_bit_number = 21;
defparam ram_block3a21.port_b_last_address = 8191;
defparam ram_block3a21.port_b_logical_ram_depth = 16384;
defparam ram_block3a21.port_b_logical_ram_width = 32;
defparam ram_block3a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_read_enable_clock = "clock1";
defparam ram_block3a21.port_b_write_enable_clock = "clock1";
defparam ram_block3a21.ram_block_type = "M9K";
defparam ram_block3a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018CF8;
// synopsys translate_on

// Location: M9K_X51_Y44_N0
cycloneive_ram_block ram_block3a54(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a54_PORTADATAOUT_bus),
	.portbdataout(ram_block3a54_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a54.clk0_core_clock_enable = "ena0";
defparam ram_block3a54.clk1_core_clock_enable = "ena1";
defparam ram_block3a54.data_interleave_offset_in_bits = 1;
defparam ram_block3a54.data_interleave_width_in_bits = 1;
defparam ram_block3a54.init_file = "meminit.hex";
defparam ram_block3a54.init_file_layout = "port_a";
defparam ram_block3a54.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a54.operation_mode = "bidir_dual_port";
defparam ram_block3a54.port_a_address_clear = "none";
defparam ram_block3a54.port_a_address_width = 13;
defparam ram_block3a54.port_a_byte_enable_clock = "none";
defparam ram_block3a54.port_a_data_out_clear = "none";
defparam ram_block3a54.port_a_data_out_clock = "none";
defparam ram_block3a54.port_a_data_width = 1;
defparam ram_block3a54.port_a_first_address = 0;
defparam ram_block3a54.port_a_first_bit_number = 22;
defparam ram_block3a54.port_a_last_address = 8191;
defparam ram_block3a54.port_a_logical_ram_depth = 16384;
defparam ram_block3a54.port_a_logical_ram_width = 32;
defparam ram_block3a54.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_address_clear = "none";
defparam ram_block3a54.port_b_address_clock = "clock1";
defparam ram_block3a54.port_b_address_width = 13;
defparam ram_block3a54.port_b_data_in_clock = "clock1";
defparam ram_block3a54.port_b_data_out_clear = "none";
defparam ram_block3a54.port_b_data_out_clock = "none";
defparam ram_block3a54.port_b_data_width = 1;
defparam ram_block3a54.port_b_first_address = 0;
defparam ram_block3a54.port_b_first_bit_number = 22;
defparam ram_block3a54.port_b_last_address = 8191;
defparam ram_block3a54.port_b_logical_ram_depth = 16384;
defparam ram_block3a54.port_b_logical_ram_width = 32;
defparam ram_block3a54.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_read_enable_clock = "clock1";
defparam ram_block3a54.port_b_write_enable_clock = "clock1";
defparam ram_block3a54.ram_block_type = "M9K";
defparam ram_block3a54.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y45_N0
cycloneive_ram_block ram_block3a22(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a22_PORTADATAOUT_bus),
	.portbdataout(ram_block3a22_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a22.clk0_core_clock_enable = "ena0";
defparam ram_block3a22.clk1_core_clock_enable = "ena1";
defparam ram_block3a22.data_interleave_offset_in_bits = 1;
defparam ram_block3a22.data_interleave_width_in_bits = 1;
defparam ram_block3a22.init_file = "meminit.hex";
defparam ram_block3a22.init_file_layout = "port_a";
defparam ram_block3a22.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a22.operation_mode = "bidir_dual_port";
defparam ram_block3a22.port_a_address_clear = "none";
defparam ram_block3a22.port_a_address_width = 13;
defparam ram_block3a22.port_a_byte_enable_clock = "none";
defparam ram_block3a22.port_a_data_out_clear = "none";
defparam ram_block3a22.port_a_data_out_clock = "none";
defparam ram_block3a22.port_a_data_width = 1;
defparam ram_block3a22.port_a_first_address = 0;
defparam ram_block3a22.port_a_first_bit_number = 22;
defparam ram_block3a22.port_a_last_address = 8191;
defparam ram_block3a22.port_a_logical_ram_depth = 16384;
defparam ram_block3a22.port_a_logical_ram_width = 32;
defparam ram_block3a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_address_clear = "none";
defparam ram_block3a22.port_b_address_clock = "clock1";
defparam ram_block3a22.port_b_address_width = 13;
defparam ram_block3a22.port_b_data_in_clock = "clock1";
defparam ram_block3a22.port_b_data_out_clear = "none";
defparam ram_block3a22.port_b_data_out_clock = "none";
defparam ram_block3a22.port_b_data_width = 1;
defparam ram_block3a22.port_b_first_address = 0;
defparam ram_block3a22.port_b_first_bit_number = 22;
defparam ram_block3a22.port_b_last_address = 8191;
defparam ram_block3a22.port_b_logical_ram_depth = 16384;
defparam ram_block3a22.port_b_logical_ram_width = 32;
defparam ram_block3a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_read_enable_clock = "clock1";
defparam ram_block3a22.port_b_write_enable_clock = "clock1";
defparam ram_block3a22.ram_block_type = "M9K";
defparam ram_block3a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010600;
// synopsys translate_on

// Location: M9K_X51_Y41_N0
cycloneive_ram_block ram_block3a55(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a55_PORTADATAOUT_bus),
	.portbdataout(ram_block3a55_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a55.clk0_core_clock_enable = "ena0";
defparam ram_block3a55.clk1_core_clock_enable = "ena1";
defparam ram_block3a55.data_interleave_offset_in_bits = 1;
defparam ram_block3a55.data_interleave_width_in_bits = 1;
defparam ram_block3a55.init_file = "meminit.hex";
defparam ram_block3a55.init_file_layout = "port_a";
defparam ram_block3a55.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a55.operation_mode = "bidir_dual_port";
defparam ram_block3a55.port_a_address_clear = "none";
defparam ram_block3a55.port_a_address_width = 13;
defparam ram_block3a55.port_a_byte_enable_clock = "none";
defparam ram_block3a55.port_a_data_out_clear = "none";
defparam ram_block3a55.port_a_data_out_clock = "none";
defparam ram_block3a55.port_a_data_width = 1;
defparam ram_block3a55.port_a_first_address = 0;
defparam ram_block3a55.port_a_first_bit_number = 23;
defparam ram_block3a55.port_a_last_address = 8191;
defparam ram_block3a55.port_a_logical_ram_depth = 16384;
defparam ram_block3a55.port_a_logical_ram_width = 32;
defparam ram_block3a55.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_address_clear = "none";
defparam ram_block3a55.port_b_address_clock = "clock1";
defparam ram_block3a55.port_b_address_width = 13;
defparam ram_block3a55.port_b_data_in_clock = "clock1";
defparam ram_block3a55.port_b_data_out_clear = "none";
defparam ram_block3a55.port_b_data_out_clock = "none";
defparam ram_block3a55.port_b_data_width = 1;
defparam ram_block3a55.port_b_first_address = 0;
defparam ram_block3a55.port_b_first_bit_number = 23;
defparam ram_block3a55.port_b_last_address = 8191;
defparam ram_block3a55.port_b_logical_ram_depth = 16384;
defparam ram_block3a55.port_b_logical_ram_width = 32;
defparam ram_block3a55.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_read_enable_clock = "clock1";
defparam ram_block3a55.port_b_write_enable_clock = "clock1";
defparam ram_block3a55.ram_block_type = "M9K";
defparam ram_block3a55.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y42_N0
cycloneive_ram_block ram_block3a23(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a23_PORTADATAOUT_bus),
	.portbdataout(ram_block3a23_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a23.clk0_core_clock_enable = "ena0";
defparam ram_block3a23.clk1_core_clock_enable = "ena1";
defparam ram_block3a23.data_interleave_offset_in_bits = 1;
defparam ram_block3a23.data_interleave_width_in_bits = 1;
defparam ram_block3a23.init_file = "meminit.hex";
defparam ram_block3a23.init_file_layout = "port_a";
defparam ram_block3a23.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a23.operation_mode = "bidir_dual_port";
defparam ram_block3a23.port_a_address_clear = "none";
defparam ram_block3a23.port_a_address_width = 13;
defparam ram_block3a23.port_a_byte_enable_clock = "none";
defparam ram_block3a23.port_a_data_out_clear = "none";
defparam ram_block3a23.port_a_data_out_clock = "none";
defparam ram_block3a23.port_a_data_width = 1;
defparam ram_block3a23.port_a_first_address = 0;
defparam ram_block3a23.port_a_first_bit_number = 23;
defparam ram_block3a23.port_a_last_address = 8191;
defparam ram_block3a23.port_a_logical_ram_depth = 16384;
defparam ram_block3a23.port_a_logical_ram_width = 32;
defparam ram_block3a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_address_clear = "none";
defparam ram_block3a23.port_b_address_clock = "clock1";
defparam ram_block3a23.port_b_address_width = 13;
defparam ram_block3a23.port_b_data_in_clock = "clock1";
defparam ram_block3a23.port_b_data_out_clear = "none";
defparam ram_block3a23.port_b_data_out_clock = "none";
defparam ram_block3a23.port_b_data_width = 1;
defparam ram_block3a23.port_b_first_address = 0;
defparam ram_block3a23.port_b_first_bit_number = 23;
defparam ram_block3a23.port_b_last_address = 8191;
defparam ram_block3a23.port_b_logical_ram_depth = 16384;
defparam ram_block3a23.port_b_logical_ram_width = 32;
defparam ram_block3a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_read_enable_clock = "clock1";
defparam ram_block3a23.port_b_write_enable_clock = "clock1";
defparam ram_block3a23.ram_block_type = "M9K";
defparam ram_block3a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001BEF8;
// synopsys translate_on

// Location: M9K_X37_Y38_N0
cycloneive_ram_block ram_block3a56(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a56_PORTADATAOUT_bus),
	.portbdataout(ram_block3a56_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a56.clk0_core_clock_enable = "ena0";
defparam ram_block3a56.clk1_core_clock_enable = "ena1";
defparam ram_block3a56.data_interleave_offset_in_bits = 1;
defparam ram_block3a56.data_interleave_width_in_bits = 1;
defparam ram_block3a56.init_file = "meminit.hex";
defparam ram_block3a56.init_file_layout = "port_a";
defparam ram_block3a56.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a56.operation_mode = "bidir_dual_port";
defparam ram_block3a56.port_a_address_clear = "none";
defparam ram_block3a56.port_a_address_width = 13;
defparam ram_block3a56.port_a_byte_enable_clock = "none";
defparam ram_block3a56.port_a_data_out_clear = "none";
defparam ram_block3a56.port_a_data_out_clock = "none";
defparam ram_block3a56.port_a_data_width = 1;
defparam ram_block3a56.port_a_first_address = 0;
defparam ram_block3a56.port_a_first_bit_number = 24;
defparam ram_block3a56.port_a_last_address = 8191;
defparam ram_block3a56.port_a_logical_ram_depth = 16384;
defparam ram_block3a56.port_a_logical_ram_width = 32;
defparam ram_block3a56.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_address_clear = "none";
defparam ram_block3a56.port_b_address_clock = "clock1";
defparam ram_block3a56.port_b_address_width = 13;
defparam ram_block3a56.port_b_data_in_clock = "clock1";
defparam ram_block3a56.port_b_data_out_clear = "none";
defparam ram_block3a56.port_b_data_out_clock = "none";
defparam ram_block3a56.port_b_data_width = 1;
defparam ram_block3a56.port_b_first_address = 0;
defparam ram_block3a56.port_b_first_bit_number = 24;
defparam ram_block3a56.port_b_last_address = 8191;
defparam ram_block3a56.port_b_logical_ram_depth = 16384;
defparam ram_block3a56.port_b_logical_ram_width = 32;
defparam ram_block3a56.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_read_enable_clock = "clock1";
defparam ram_block3a56.port_b_write_enable_clock = "clock1";
defparam ram_block3a56.ram_block_type = "M9K";
defparam ram_block3a56.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y35_N0
cycloneive_ram_block ram_block3a24(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a24_PORTADATAOUT_bus),
	.portbdataout(ram_block3a24_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a24.clk0_core_clock_enable = "ena0";
defparam ram_block3a24.clk1_core_clock_enable = "ena1";
defparam ram_block3a24.data_interleave_offset_in_bits = 1;
defparam ram_block3a24.data_interleave_width_in_bits = 1;
defparam ram_block3a24.init_file = "meminit.hex";
defparam ram_block3a24.init_file_layout = "port_a";
defparam ram_block3a24.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a24.operation_mode = "bidir_dual_port";
defparam ram_block3a24.port_a_address_clear = "none";
defparam ram_block3a24.port_a_address_width = 13;
defparam ram_block3a24.port_a_byte_enable_clock = "none";
defparam ram_block3a24.port_a_data_out_clear = "none";
defparam ram_block3a24.port_a_data_out_clock = "none";
defparam ram_block3a24.port_a_data_width = 1;
defparam ram_block3a24.port_a_first_address = 0;
defparam ram_block3a24.port_a_first_bit_number = 24;
defparam ram_block3a24.port_a_last_address = 8191;
defparam ram_block3a24.port_a_logical_ram_depth = 16384;
defparam ram_block3a24.port_a_logical_ram_width = 32;
defparam ram_block3a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_address_clear = "none";
defparam ram_block3a24.port_b_address_clock = "clock1";
defparam ram_block3a24.port_b_address_width = 13;
defparam ram_block3a24.port_b_data_in_clock = "clock1";
defparam ram_block3a24.port_b_data_out_clear = "none";
defparam ram_block3a24.port_b_data_out_clock = "none";
defparam ram_block3a24.port_b_data_width = 1;
defparam ram_block3a24.port_b_first_address = 0;
defparam ram_block3a24.port_b_first_bit_number = 24;
defparam ram_block3a24.port_b_last_address = 8191;
defparam ram_block3a24.port_b_logical_ram_depth = 16384;
defparam ram_block3a24.port_b_logical_ram_width = 32;
defparam ram_block3a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_read_enable_clock = "clock1";
defparam ram_block3a24.port_b_write_enable_clock = "clock1";
defparam ram_block3a24.ram_block_type = "M9K";
defparam ram_block3a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018078;
// synopsys translate_on

// Location: M9K_X51_Y38_N0
cycloneive_ram_block ram_block3a57(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a57_PORTADATAOUT_bus),
	.portbdataout(ram_block3a57_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a57.clk0_core_clock_enable = "ena0";
defparam ram_block3a57.clk1_core_clock_enable = "ena1";
defparam ram_block3a57.data_interleave_offset_in_bits = 1;
defparam ram_block3a57.data_interleave_width_in_bits = 1;
defparam ram_block3a57.init_file = "meminit.hex";
defparam ram_block3a57.init_file_layout = "port_a";
defparam ram_block3a57.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a57.operation_mode = "bidir_dual_port";
defparam ram_block3a57.port_a_address_clear = "none";
defparam ram_block3a57.port_a_address_width = 13;
defparam ram_block3a57.port_a_byte_enable_clock = "none";
defparam ram_block3a57.port_a_data_out_clear = "none";
defparam ram_block3a57.port_a_data_out_clock = "none";
defparam ram_block3a57.port_a_data_width = 1;
defparam ram_block3a57.port_a_first_address = 0;
defparam ram_block3a57.port_a_first_bit_number = 25;
defparam ram_block3a57.port_a_last_address = 8191;
defparam ram_block3a57.port_a_logical_ram_depth = 16384;
defparam ram_block3a57.port_a_logical_ram_width = 32;
defparam ram_block3a57.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_address_clear = "none";
defparam ram_block3a57.port_b_address_clock = "clock1";
defparam ram_block3a57.port_b_address_width = 13;
defparam ram_block3a57.port_b_data_in_clock = "clock1";
defparam ram_block3a57.port_b_data_out_clear = "none";
defparam ram_block3a57.port_b_data_out_clock = "none";
defparam ram_block3a57.port_b_data_width = 1;
defparam ram_block3a57.port_b_first_address = 0;
defparam ram_block3a57.port_b_first_bit_number = 25;
defparam ram_block3a57.port_b_last_address = 8191;
defparam ram_block3a57.port_b_logical_ram_depth = 16384;
defparam ram_block3a57.port_b_logical_ram_width = 32;
defparam ram_block3a57.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_read_enable_clock = "clock1";
defparam ram_block3a57.port_b_write_enable_clock = "clock1";
defparam ram_block3a57.ram_block_type = "M9K";
defparam ram_block3a57.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y37_N0
cycloneive_ram_block ram_block3a25(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a25_PORTADATAOUT_bus),
	.portbdataout(ram_block3a25_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a25.clk0_core_clock_enable = "ena0";
defparam ram_block3a25.clk1_core_clock_enable = "ena1";
defparam ram_block3a25.data_interleave_offset_in_bits = 1;
defparam ram_block3a25.data_interleave_width_in_bits = 1;
defparam ram_block3a25.init_file = "meminit.hex";
defparam ram_block3a25.init_file_layout = "port_a";
defparam ram_block3a25.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a25.operation_mode = "bidir_dual_port";
defparam ram_block3a25.port_a_address_clear = "none";
defparam ram_block3a25.port_a_address_width = 13;
defparam ram_block3a25.port_a_byte_enable_clock = "none";
defparam ram_block3a25.port_a_data_out_clear = "none";
defparam ram_block3a25.port_a_data_out_clock = "none";
defparam ram_block3a25.port_a_data_width = 1;
defparam ram_block3a25.port_a_first_address = 0;
defparam ram_block3a25.port_a_first_bit_number = 25;
defparam ram_block3a25.port_a_last_address = 8191;
defparam ram_block3a25.port_a_logical_ram_depth = 16384;
defparam ram_block3a25.port_a_logical_ram_width = 32;
defparam ram_block3a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_address_clear = "none";
defparam ram_block3a25.port_b_address_clock = "clock1";
defparam ram_block3a25.port_b_address_width = 13;
defparam ram_block3a25.port_b_data_in_clock = "clock1";
defparam ram_block3a25.port_b_data_out_clear = "none";
defparam ram_block3a25.port_b_data_out_clock = "none";
defparam ram_block3a25.port_b_data_width = 1;
defparam ram_block3a25.port_b_first_address = 0;
defparam ram_block3a25.port_b_first_bit_number = 25;
defparam ram_block3a25.port_b_last_address = 8191;
defparam ram_block3a25.port_b_logical_ram_depth = 16384;
defparam ram_block3a25.port_b_logical_ram_width = 32;
defparam ram_block3a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_read_enable_clock = "clock1";
defparam ram_block3a25.port_b_write_enable_clock = "clock1";
defparam ram_block3a25.ram_block_type = "M9K";
defparam ram_block3a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018078;
// synopsys translate_on

// Location: M9K_X37_Y42_N0
cycloneive_ram_block ram_block3a58(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a58_PORTADATAOUT_bus),
	.portbdataout(ram_block3a58_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a58.clk0_core_clock_enable = "ena0";
defparam ram_block3a58.clk1_core_clock_enable = "ena1";
defparam ram_block3a58.data_interleave_offset_in_bits = 1;
defparam ram_block3a58.data_interleave_width_in_bits = 1;
defparam ram_block3a58.init_file = "meminit.hex";
defparam ram_block3a58.init_file_layout = "port_a";
defparam ram_block3a58.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a58.operation_mode = "bidir_dual_port";
defparam ram_block3a58.port_a_address_clear = "none";
defparam ram_block3a58.port_a_address_width = 13;
defparam ram_block3a58.port_a_byte_enable_clock = "none";
defparam ram_block3a58.port_a_data_out_clear = "none";
defparam ram_block3a58.port_a_data_out_clock = "none";
defparam ram_block3a58.port_a_data_width = 1;
defparam ram_block3a58.port_a_first_address = 0;
defparam ram_block3a58.port_a_first_bit_number = 26;
defparam ram_block3a58.port_a_last_address = 8191;
defparam ram_block3a58.port_a_logical_ram_depth = 16384;
defparam ram_block3a58.port_a_logical_ram_width = 32;
defparam ram_block3a58.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_address_clear = "none";
defparam ram_block3a58.port_b_address_clock = "clock1";
defparam ram_block3a58.port_b_address_width = 13;
defparam ram_block3a58.port_b_data_in_clock = "clock1";
defparam ram_block3a58.port_b_data_out_clear = "none";
defparam ram_block3a58.port_b_data_out_clock = "none";
defparam ram_block3a58.port_b_data_width = 1;
defparam ram_block3a58.port_b_first_address = 0;
defparam ram_block3a58.port_b_first_bit_number = 26;
defparam ram_block3a58.port_b_last_address = 8191;
defparam ram_block3a58.port_b_logical_ram_depth = 16384;
defparam ram_block3a58.port_b_logical_ram_width = 32;
defparam ram_block3a58.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_read_enable_clock = "clock1";
defparam ram_block3a58.port_b_write_enable_clock = "clock1";
defparam ram_block3a58.ram_block_type = "M9K";
defparam ram_block3a58.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y41_N0
cycloneive_ram_block ram_block3a26(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a26_PORTADATAOUT_bus),
	.portbdataout(ram_block3a26_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a26.clk0_core_clock_enable = "ena0";
defparam ram_block3a26.clk1_core_clock_enable = "ena1";
defparam ram_block3a26.data_interleave_offset_in_bits = 1;
defparam ram_block3a26.data_interleave_width_in_bits = 1;
defparam ram_block3a26.init_file = "meminit.hex";
defparam ram_block3a26.init_file_layout = "port_a";
defparam ram_block3a26.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a26.operation_mode = "bidir_dual_port";
defparam ram_block3a26.port_a_address_clear = "none";
defparam ram_block3a26.port_a_address_width = 13;
defparam ram_block3a26.port_a_byte_enable_clock = "none";
defparam ram_block3a26.port_a_data_out_clear = "none";
defparam ram_block3a26.port_a_data_out_clock = "none";
defparam ram_block3a26.port_a_data_width = 1;
defparam ram_block3a26.port_a_first_address = 0;
defparam ram_block3a26.port_a_first_bit_number = 26;
defparam ram_block3a26.port_a_last_address = 8191;
defparam ram_block3a26.port_a_logical_ram_depth = 16384;
defparam ram_block3a26.port_a_logical_ram_width = 32;
defparam ram_block3a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_address_clear = "none";
defparam ram_block3a26.port_b_address_clock = "clock1";
defparam ram_block3a26.port_b_address_width = 13;
defparam ram_block3a26.port_b_data_in_clock = "clock1";
defparam ram_block3a26.port_b_data_out_clear = "none";
defparam ram_block3a26.port_b_data_out_clock = "none";
defparam ram_block3a26.port_b_data_width = 1;
defparam ram_block3a26.port_b_first_address = 0;
defparam ram_block3a26.port_b_first_bit_number = 26;
defparam ram_block3a26.port_b_last_address = 8191;
defparam ram_block3a26.port_b_logical_ram_depth = 16384;
defparam ram_block3a26.port_b_logical_ram_width = 32;
defparam ram_block3a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_read_enable_clock = "clock1";
defparam ram_block3a26.port_b_write_enable_clock = "clock1";
defparam ram_block3a26.ram_block_type = "M9K";
defparam ram_block3a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000180FF;
// synopsys translate_on

// Location: M9K_X37_Y45_N0
cycloneive_ram_block ram_block3a59(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a59_PORTADATAOUT_bus),
	.portbdataout(ram_block3a59_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a59.clk0_core_clock_enable = "ena0";
defparam ram_block3a59.clk1_core_clock_enable = "ena1";
defparam ram_block3a59.data_interleave_offset_in_bits = 1;
defparam ram_block3a59.data_interleave_width_in_bits = 1;
defparam ram_block3a59.init_file = "meminit.hex";
defparam ram_block3a59.init_file_layout = "port_a";
defparam ram_block3a59.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a59.operation_mode = "bidir_dual_port";
defparam ram_block3a59.port_a_address_clear = "none";
defparam ram_block3a59.port_a_address_width = 13;
defparam ram_block3a59.port_a_byte_enable_clock = "none";
defparam ram_block3a59.port_a_data_out_clear = "none";
defparam ram_block3a59.port_a_data_out_clock = "none";
defparam ram_block3a59.port_a_data_width = 1;
defparam ram_block3a59.port_a_first_address = 0;
defparam ram_block3a59.port_a_first_bit_number = 27;
defparam ram_block3a59.port_a_last_address = 8191;
defparam ram_block3a59.port_a_logical_ram_depth = 16384;
defparam ram_block3a59.port_a_logical_ram_width = 32;
defparam ram_block3a59.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_address_clear = "none";
defparam ram_block3a59.port_b_address_clock = "clock1";
defparam ram_block3a59.port_b_address_width = 13;
defparam ram_block3a59.port_b_data_in_clock = "clock1";
defparam ram_block3a59.port_b_data_out_clear = "none";
defparam ram_block3a59.port_b_data_out_clock = "none";
defparam ram_block3a59.port_b_data_width = 1;
defparam ram_block3a59.port_b_first_address = 0;
defparam ram_block3a59.port_b_first_bit_number = 27;
defparam ram_block3a59.port_b_last_address = 8191;
defparam ram_block3a59.port_b_logical_ram_depth = 16384;
defparam ram_block3a59.port_b_logical_ram_width = 32;
defparam ram_block3a59.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_read_enable_clock = "clock1";
defparam ram_block3a59.port_b_write_enable_clock = "clock1";
defparam ram_block3a59.ram_block_type = "M9K";
defparam ram_block3a59.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y45_N0
cycloneive_ram_block ram_block3a27(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a27_PORTADATAOUT_bus),
	.portbdataout(ram_block3a27_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a27.clk0_core_clock_enable = "ena0";
defparam ram_block3a27.clk1_core_clock_enable = "ena1";
defparam ram_block3a27.data_interleave_offset_in_bits = 1;
defparam ram_block3a27.data_interleave_width_in_bits = 1;
defparam ram_block3a27.init_file = "meminit.hex";
defparam ram_block3a27.init_file_layout = "port_a";
defparam ram_block3a27.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a27.operation_mode = "bidir_dual_port";
defparam ram_block3a27.port_a_address_clear = "none";
defparam ram_block3a27.port_a_address_width = 13;
defparam ram_block3a27.port_a_byte_enable_clock = "none";
defparam ram_block3a27.port_a_data_out_clear = "none";
defparam ram_block3a27.port_a_data_out_clock = "none";
defparam ram_block3a27.port_a_data_width = 1;
defparam ram_block3a27.port_a_first_address = 0;
defparam ram_block3a27.port_a_first_bit_number = 27;
defparam ram_block3a27.port_a_last_address = 8191;
defparam ram_block3a27.port_a_logical_ram_depth = 16384;
defparam ram_block3a27.port_a_logical_ram_width = 32;
defparam ram_block3a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_address_clear = "none";
defparam ram_block3a27.port_b_address_clock = "clock1";
defparam ram_block3a27.port_b_address_width = 13;
defparam ram_block3a27.port_b_data_in_clock = "clock1";
defparam ram_block3a27.port_b_data_out_clear = "none";
defparam ram_block3a27.port_b_data_out_clock = "none";
defparam ram_block3a27.port_b_data_width = 1;
defparam ram_block3a27.port_b_first_address = 0;
defparam ram_block3a27.port_b_first_bit_number = 27;
defparam ram_block3a27.port_b_last_address = 8191;
defparam ram_block3a27.port_b_logical_ram_depth = 16384;
defparam ram_block3a27.port_b_logical_ram_width = 32;
defparam ram_block3a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_read_enable_clock = "clock1";
defparam ram_block3a27.port_b_write_enable_clock = "clock1";
defparam ram_block3a27.ram_block_type = "M9K";
defparam ram_block3a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000180B8;
// synopsys translate_on

// Location: M9K_X64_Y36_N0
cycloneive_ram_block ram_block3a60(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a60_PORTADATAOUT_bus),
	.portbdataout(ram_block3a60_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a60.clk0_core_clock_enable = "ena0";
defparam ram_block3a60.clk1_core_clock_enable = "ena1";
defparam ram_block3a60.data_interleave_offset_in_bits = 1;
defparam ram_block3a60.data_interleave_width_in_bits = 1;
defparam ram_block3a60.init_file = "meminit.hex";
defparam ram_block3a60.init_file_layout = "port_a";
defparam ram_block3a60.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a60.operation_mode = "bidir_dual_port";
defparam ram_block3a60.port_a_address_clear = "none";
defparam ram_block3a60.port_a_address_width = 13;
defparam ram_block3a60.port_a_byte_enable_clock = "none";
defparam ram_block3a60.port_a_data_out_clear = "none";
defparam ram_block3a60.port_a_data_out_clock = "none";
defparam ram_block3a60.port_a_data_width = 1;
defparam ram_block3a60.port_a_first_address = 0;
defparam ram_block3a60.port_a_first_bit_number = 28;
defparam ram_block3a60.port_a_last_address = 8191;
defparam ram_block3a60.port_a_logical_ram_depth = 16384;
defparam ram_block3a60.port_a_logical_ram_width = 32;
defparam ram_block3a60.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_address_clear = "none";
defparam ram_block3a60.port_b_address_clock = "clock1";
defparam ram_block3a60.port_b_address_width = 13;
defparam ram_block3a60.port_b_data_in_clock = "clock1";
defparam ram_block3a60.port_b_data_out_clear = "none";
defparam ram_block3a60.port_b_data_out_clock = "none";
defparam ram_block3a60.port_b_data_width = 1;
defparam ram_block3a60.port_b_first_address = 0;
defparam ram_block3a60.port_b_first_bit_number = 28;
defparam ram_block3a60.port_b_last_address = 8191;
defparam ram_block3a60.port_b_logical_ram_depth = 16384;
defparam ram_block3a60.port_b_logical_ram_width = 32;
defparam ram_block3a60.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_read_enable_clock = "clock1";
defparam ram_block3a60.port_b_write_enable_clock = "clock1";
defparam ram_block3a60.ram_block_type = "M9K";
defparam ram_block3a60.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y36_N0
cycloneive_ram_block ram_block3a28(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a28_PORTADATAOUT_bus),
	.portbdataout(ram_block3a28_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a28.clk0_core_clock_enable = "ena0";
defparam ram_block3a28.clk1_core_clock_enable = "ena1";
defparam ram_block3a28.data_interleave_offset_in_bits = 1;
defparam ram_block3a28.data_interleave_width_in_bits = 1;
defparam ram_block3a28.init_file = "meminit.hex";
defparam ram_block3a28.init_file_layout = "port_a";
defparam ram_block3a28.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a28.operation_mode = "bidir_dual_port";
defparam ram_block3a28.port_a_address_clear = "none";
defparam ram_block3a28.port_a_address_width = 13;
defparam ram_block3a28.port_a_byte_enable_clock = "none";
defparam ram_block3a28.port_a_data_out_clear = "none";
defparam ram_block3a28.port_a_data_out_clock = "none";
defparam ram_block3a28.port_a_data_width = 1;
defparam ram_block3a28.port_a_first_address = 0;
defparam ram_block3a28.port_a_first_bit_number = 28;
defparam ram_block3a28.port_a_last_address = 8191;
defparam ram_block3a28.port_a_logical_ram_depth = 16384;
defparam ram_block3a28.port_a_logical_ram_width = 32;
defparam ram_block3a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_address_clear = "none";
defparam ram_block3a28.port_b_address_clock = "clock1";
defparam ram_block3a28.port_b_address_width = 13;
defparam ram_block3a28.port_b_data_in_clock = "clock1";
defparam ram_block3a28.port_b_data_out_clear = "none";
defparam ram_block3a28.port_b_data_out_clock = "none";
defparam ram_block3a28.port_b_data_width = 1;
defparam ram_block3a28.port_b_first_address = 0;
defparam ram_block3a28.port_b_first_bit_number = 28;
defparam ram_block3a28.port_b_last_address = 8191;
defparam ram_block3a28.port_b_logical_ram_depth = 16384;
defparam ram_block3a28.port_b_logical_ram_width = 32;
defparam ram_block3a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_read_enable_clock = "clock1";
defparam ram_block3a28.port_b_write_enable_clock = "clock1";
defparam ram_block3a28.ram_block_type = "M9K";
defparam ram_block3a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000016407;
// synopsys translate_on

// Location: M9K_X51_Y32_N0
cycloneive_ram_block ram_block3a61(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a61_PORTADATAOUT_bus),
	.portbdataout(ram_block3a61_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a61.clk0_core_clock_enable = "ena0";
defparam ram_block3a61.clk1_core_clock_enable = "ena1";
defparam ram_block3a61.data_interleave_offset_in_bits = 1;
defparam ram_block3a61.data_interleave_width_in_bits = 1;
defparam ram_block3a61.init_file = "meminit.hex";
defparam ram_block3a61.init_file_layout = "port_a";
defparam ram_block3a61.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a61.operation_mode = "bidir_dual_port";
defparam ram_block3a61.port_a_address_clear = "none";
defparam ram_block3a61.port_a_address_width = 13;
defparam ram_block3a61.port_a_byte_enable_clock = "none";
defparam ram_block3a61.port_a_data_out_clear = "none";
defparam ram_block3a61.port_a_data_out_clock = "none";
defparam ram_block3a61.port_a_data_width = 1;
defparam ram_block3a61.port_a_first_address = 0;
defparam ram_block3a61.port_a_first_bit_number = 29;
defparam ram_block3a61.port_a_last_address = 8191;
defparam ram_block3a61.port_a_logical_ram_depth = 16384;
defparam ram_block3a61.port_a_logical_ram_width = 32;
defparam ram_block3a61.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_address_clear = "none";
defparam ram_block3a61.port_b_address_clock = "clock1";
defparam ram_block3a61.port_b_address_width = 13;
defparam ram_block3a61.port_b_data_in_clock = "clock1";
defparam ram_block3a61.port_b_data_out_clear = "none";
defparam ram_block3a61.port_b_data_out_clock = "none";
defparam ram_block3a61.port_b_data_width = 1;
defparam ram_block3a61.port_b_first_address = 0;
defparam ram_block3a61.port_b_first_bit_number = 29;
defparam ram_block3a61.port_b_last_address = 8191;
defparam ram_block3a61.port_b_logical_ram_depth = 16384;
defparam ram_block3a61.port_b_logical_ram_width = 32;
defparam ram_block3a61.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_read_enable_clock = "clock1";
defparam ram_block3a61.port_b_write_enable_clock = "clock1";
defparam ram_block3a61.ram_block_type = "M9K";
defparam ram_block3a61.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y33_N0
cycloneive_ram_block ram_block3a29(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a29_PORTADATAOUT_bus),
	.portbdataout(ram_block3a29_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a29.clk0_core_clock_enable = "ena0";
defparam ram_block3a29.clk1_core_clock_enable = "ena1";
defparam ram_block3a29.data_interleave_offset_in_bits = 1;
defparam ram_block3a29.data_interleave_width_in_bits = 1;
defparam ram_block3a29.init_file = "meminit.hex";
defparam ram_block3a29.init_file_layout = "port_a";
defparam ram_block3a29.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a29.operation_mode = "bidir_dual_port";
defparam ram_block3a29.port_a_address_clear = "none";
defparam ram_block3a29.port_a_address_width = 13;
defparam ram_block3a29.port_a_byte_enable_clock = "none";
defparam ram_block3a29.port_a_data_out_clear = "none";
defparam ram_block3a29.port_a_data_out_clock = "none";
defparam ram_block3a29.port_a_data_width = 1;
defparam ram_block3a29.port_a_first_address = 0;
defparam ram_block3a29.port_a_first_bit_number = 29;
defparam ram_block3a29.port_a_last_address = 8191;
defparam ram_block3a29.port_a_logical_ram_depth = 16384;
defparam ram_block3a29.port_a_logical_ram_width = 32;
defparam ram_block3a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_address_clear = "none";
defparam ram_block3a29.port_b_address_clock = "clock1";
defparam ram_block3a29.port_b_address_width = 13;
defparam ram_block3a29.port_b_data_in_clock = "clock1";
defparam ram_block3a29.port_b_data_out_clear = "none";
defparam ram_block3a29.port_b_data_out_clock = "none";
defparam ram_block3a29.port_b_data_width = 1;
defparam ram_block3a29.port_b_first_address = 0;
defparam ram_block3a29.port_b_first_bit_number = 29;
defparam ram_block3a29.port_b_last_address = 8191;
defparam ram_block3a29.port_b_logical_ram_depth = 16384;
defparam ram_block3a29.port_b_logical_ram_width = 32;
defparam ram_block3a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_read_enable_clock = "clock1";
defparam ram_block3a29.port_b_write_enable_clock = "clock1";
defparam ram_block3a29.ram_block_type = "M9K";
defparam ram_block3a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001804F;
// synopsys translate_on

// Location: M9K_X64_Y38_N0
cycloneive_ram_block ram_block3a62(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a62_PORTADATAOUT_bus),
	.portbdataout(ram_block3a62_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a62.clk0_core_clock_enable = "ena0";
defparam ram_block3a62.clk1_core_clock_enable = "ena1";
defparam ram_block3a62.data_interleave_offset_in_bits = 1;
defparam ram_block3a62.data_interleave_width_in_bits = 1;
defparam ram_block3a62.init_file = "meminit.hex";
defparam ram_block3a62.init_file_layout = "port_a";
defparam ram_block3a62.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a62.operation_mode = "bidir_dual_port";
defparam ram_block3a62.port_a_address_clear = "none";
defparam ram_block3a62.port_a_address_width = 13;
defparam ram_block3a62.port_a_byte_enable_clock = "none";
defparam ram_block3a62.port_a_data_out_clear = "none";
defparam ram_block3a62.port_a_data_out_clock = "none";
defparam ram_block3a62.port_a_data_width = 1;
defparam ram_block3a62.port_a_first_address = 0;
defparam ram_block3a62.port_a_first_bit_number = 30;
defparam ram_block3a62.port_a_last_address = 8191;
defparam ram_block3a62.port_a_logical_ram_depth = 16384;
defparam ram_block3a62.port_a_logical_ram_width = 32;
defparam ram_block3a62.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_address_clear = "none";
defparam ram_block3a62.port_b_address_clock = "clock1";
defparam ram_block3a62.port_b_address_width = 13;
defparam ram_block3a62.port_b_data_in_clock = "clock1";
defparam ram_block3a62.port_b_data_out_clear = "none";
defparam ram_block3a62.port_b_data_out_clock = "none";
defparam ram_block3a62.port_b_data_width = 1;
defparam ram_block3a62.port_b_first_address = 0;
defparam ram_block3a62.port_b_first_bit_number = 30;
defparam ram_block3a62.port_b_last_address = 8191;
defparam ram_block3a62.port_b_logical_ram_depth = 16384;
defparam ram_block3a62.port_b_logical_ram_width = 32;
defparam ram_block3a62.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_read_enable_clock = "clock1";
defparam ram_block3a62.port_b_write_enable_clock = "clock1";
defparam ram_block3a62.ram_block_type = "M9K";
defparam ram_block3a62.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y37_N0
cycloneive_ram_block ram_block3a30(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a30_PORTADATAOUT_bus),
	.portbdataout(ram_block3a30_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a30.clk0_core_clock_enable = "ena0";
defparam ram_block3a30.clk1_core_clock_enable = "ena1";
defparam ram_block3a30.data_interleave_offset_in_bits = 1;
defparam ram_block3a30.data_interleave_width_in_bits = 1;
defparam ram_block3a30.init_file = "meminit.hex";
defparam ram_block3a30.init_file_layout = "port_a";
defparam ram_block3a30.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a30.operation_mode = "bidir_dual_port";
defparam ram_block3a30.port_a_address_clear = "none";
defparam ram_block3a30.port_a_address_width = 13;
defparam ram_block3a30.port_a_byte_enable_clock = "none";
defparam ram_block3a30.port_a_data_out_clear = "none";
defparam ram_block3a30.port_a_data_out_clock = "none";
defparam ram_block3a30.port_a_data_width = 1;
defparam ram_block3a30.port_a_first_address = 0;
defparam ram_block3a30.port_a_first_bit_number = 30;
defparam ram_block3a30.port_a_last_address = 8191;
defparam ram_block3a30.port_a_logical_ram_depth = 16384;
defparam ram_block3a30.port_a_logical_ram_width = 32;
defparam ram_block3a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_address_clear = "none";
defparam ram_block3a30.port_b_address_clock = "clock1";
defparam ram_block3a30.port_b_address_width = 13;
defparam ram_block3a30.port_b_data_in_clock = "clock1";
defparam ram_block3a30.port_b_data_out_clear = "none";
defparam ram_block3a30.port_b_data_out_clock = "none";
defparam ram_block3a30.port_b_data_width = 1;
defparam ram_block3a30.port_b_first_address = 0;
defparam ram_block3a30.port_b_first_bit_number = 30;
defparam ram_block3a30.port_b_last_address = 8191;
defparam ram_block3a30.port_b_logical_ram_depth = 16384;
defparam ram_block3a30.port_b_logical_ram_width = 32;
defparam ram_block3a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_read_enable_clock = "clock1";
defparam ram_block3a30.port_b_write_enable_clock = "clock1";
defparam ram_block3a30.ram_block_type = "M9K";
defparam ram_block3a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
// synopsys translate_on

// Location: M9K_X37_Y40_N0
cycloneive_ram_block ram_block3a63(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a63_PORTADATAOUT_bus),
	.portbdataout(ram_block3a63_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a63.clk0_core_clock_enable = "ena0";
defparam ram_block3a63.clk1_core_clock_enable = "ena1";
defparam ram_block3a63.data_interleave_offset_in_bits = 1;
defparam ram_block3a63.data_interleave_width_in_bits = 1;
defparam ram_block3a63.init_file = "meminit.hex";
defparam ram_block3a63.init_file_layout = "port_a";
defparam ram_block3a63.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a63.operation_mode = "bidir_dual_port";
defparam ram_block3a63.port_a_address_clear = "none";
defparam ram_block3a63.port_a_address_width = 13;
defparam ram_block3a63.port_a_byte_enable_clock = "none";
defparam ram_block3a63.port_a_data_out_clear = "none";
defparam ram_block3a63.port_a_data_out_clock = "none";
defparam ram_block3a63.port_a_data_width = 1;
defparam ram_block3a63.port_a_first_address = 0;
defparam ram_block3a63.port_a_first_bit_number = 31;
defparam ram_block3a63.port_a_last_address = 8191;
defparam ram_block3a63.port_a_logical_ram_depth = 16384;
defparam ram_block3a63.port_a_logical_ram_width = 32;
defparam ram_block3a63.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_address_clear = "none";
defparam ram_block3a63.port_b_address_clock = "clock1";
defparam ram_block3a63.port_b_address_width = 13;
defparam ram_block3a63.port_b_data_in_clock = "clock1";
defparam ram_block3a63.port_b_data_out_clear = "none";
defparam ram_block3a63.port_b_data_out_clock = "none";
defparam ram_block3a63.port_b_data_width = 1;
defparam ram_block3a63.port_b_first_address = 0;
defparam ram_block3a63.port_b_first_bit_number = 31;
defparam ram_block3a63.port_b_last_address = 8191;
defparam ram_block3a63.port_b_logical_ram_depth = 16384;
defparam ram_block3a63.port_b_logical_ram_width = 32;
defparam ram_block3a63.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_read_enable_clock = "clock1";
defparam ram_block3a63.port_b_write_enable_clock = "clock1";
defparam ram_block3a63.ram_block_type = "M9K";
defparam ram_block3a63.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y40_N0
cycloneive_ram_block ram_block3a31(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a31_PORTADATAOUT_bus),
	.portbdataout(ram_block3a31_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a31.clk0_core_clock_enable = "ena0";
defparam ram_block3a31.clk1_core_clock_enable = "ena1";
defparam ram_block3a31.data_interleave_offset_in_bits = 1;
defparam ram_block3a31.data_interleave_width_in_bits = 1;
defparam ram_block3a31.init_file = "meminit.hex";
defparam ram_block3a31.init_file_layout = "port_a";
defparam ram_block3a31.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a31.operation_mode = "bidir_dual_port";
defparam ram_block3a31.port_a_address_clear = "none";
defparam ram_block3a31.port_a_address_width = 13;
defparam ram_block3a31.port_a_byte_enable_clock = "none";
defparam ram_block3a31.port_a_data_out_clear = "none";
defparam ram_block3a31.port_a_data_out_clock = "none";
defparam ram_block3a31.port_a_data_width = 1;
defparam ram_block3a31.port_a_first_address = 0;
defparam ram_block3a31.port_a_first_bit_number = 31;
defparam ram_block3a31.port_a_last_address = 8191;
defparam ram_block3a31.port_a_logical_ram_depth = 16384;
defparam ram_block3a31.port_a_logical_ram_width = 32;
defparam ram_block3a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_address_clear = "none";
defparam ram_block3a31.port_b_address_clock = "clock1";
defparam ram_block3a31.port_b_address_width = 13;
defparam ram_block3a31.port_b_data_in_clock = "clock1";
defparam ram_block3a31.port_b_data_out_clear = "none";
defparam ram_block3a31.port_b_data_out_clock = "none";
defparam ram_block3a31.port_b_data_width = 1;
defparam ram_block3a31.port_b_first_address = 0;
defparam ram_block3a31.port_b_first_bit_number = 31;
defparam ram_block3a31.port_b_last_address = 8191;
defparam ram_block3a31.port_b_logical_ram_depth = 16384;
defparam ram_block3a31.port_b_logical_ram_width = 32;
defparam ram_block3a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_read_enable_clock = "clock1";
defparam ram_block3a31.port_b_write_enable_clock = "clock1";
defparam ram_block3a31.ram_block_type = "M9K";
defparam ram_block3a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000180B8;
// synopsys translate_on

// Location: FF_X66_Y38_N31
dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(gnd),
	.asdata(ramaddr1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_a_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N19
dffeas \address_reg_b[0] (
	.clk(clock1),
	.d(\address_reg_b[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_b_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_b[0] .is_wysiwyg = "true";
defparam \address_reg_b[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N18
cycloneive_lcell_comb \address_reg_b[0]~feeder (
// Equation(s):
// \address_reg_b[0]~feeder_combout  = ram_rom_addr_reg_13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_13),
	.cin(gnd),
	.combout(\address_reg_b[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \address_reg_b[0]~feeder .lut_mask = 16'hFF00;
defparam \address_reg_b[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa (
	ramaddr,
	always1,
	ramWEN,
	eq_node_1,
	eq_node_0,
	devpor,
	devclrn,
	devoe);
input 	ramaddr;
input 	always1;
input 	ramWEN;
output 	eq_node_1;
output 	eq_node_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X61_Y40_N8
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (always1 & (\ramWEN~0_combout  & !\ramaddr~25_combout ))

	.dataa(always1),
	.datab(gnd),
	.datac(ramWEN),
	.datad(ramaddr),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h00A0;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N0
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (always1 & (\ramWEN~0_combout  & \ramaddr~25_combout ))

	.dataa(always1),
	.datab(gnd),
	.datac(ramWEN),
	.datad(ramaddr),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'hA000;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa_1 (
	ram_rom_addr_reg_13,
	sdr,
	eq_node_1,
	eq_node_0,
	irf_reg_2_1,
	state_5,
	devpor,
	devclrn,
	devoe);
input 	ram_rom_addr_reg_13;
input 	sdr;
output 	eq_node_1;
output 	eq_node_0;
input 	irf_reg_2_1;
input 	state_5;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X45_Y39_N14
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & (ram_rom_addr_reg_13 & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & sdr)))

	.dataa(irf_reg_2_1),
	.datab(ram_rom_addr_reg_13),
	.datac(state_5),
	.datad(sdr),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h8000;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N28
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & (!ram_rom_addr_reg_13 & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & sdr)))

	.dataa(irf_reg_2_1),
	.datab(ram_rom_addr_reg_13),
	.datac(state_5),
	.datad(sdr),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h2000;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_mod_ram_rom (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg1,
	ram_rom_data_reg_0,
	ram_rom_addr_reg_13,
	ram_rom_addr_reg_0,
	ram_rom_addr_reg_1,
	ram_rom_addr_reg_2,
	ram_rom_addr_reg_3,
	ram_rom_addr_reg_4,
	ram_rom_addr_reg_5,
	ram_rom_addr_reg_6,
	ram_rom_addr_reg_7,
	ram_rom_addr_reg_8,
	ram_rom_addr_reg_9,
	ram_rom_addr_reg_10,
	ram_rom_addr_reg_11,
	ram_rom_addr_reg_12,
	ram_rom_data_reg_1,
	ram_rom_data_reg_2,
	ram_rom_data_reg_3,
	ram_rom_data_reg_4,
	ram_rom_data_reg_5,
	ram_rom_data_reg_6,
	ram_rom_data_reg_7,
	ram_rom_data_reg_8,
	ram_rom_data_reg_9,
	ram_rom_data_reg_10,
	ram_rom_data_reg_11,
	ram_rom_data_reg_12,
	ram_rom_data_reg_13,
	ram_rom_data_reg_14,
	ram_rom_data_reg_15,
	ram_rom_data_reg_16,
	ram_rom_data_reg_17,
	ram_rom_data_reg_18,
	ram_rom_data_reg_19,
	ram_rom_data_reg_20,
	ram_rom_data_reg_21,
	ram_rom_data_reg_22,
	ram_rom_data_reg_23,
	ram_rom_data_reg_24,
	ram_rom_data_reg_25,
	ram_rom_data_reg_26,
	ram_rom_data_reg_27,
	ram_rom_data_reg_28,
	ram_rom_data_reg_29,
	ram_rom_data_reg_30,
	ram_rom_data_reg_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	sdr,
	address_reg_b_0,
	altera_internal_jtag,
	state_4,
	ir_in,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_4_1,
	node_ena_1,
	clr,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	raw_tck,
	devpor,
	devclrn,
	devoe);
input 	ram_block3a32;
input 	ram_block3a0;
input 	ram_block3a33;
input 	ram_block3a1;
input 	ram_block3a34;
input 	ram_block3a2;
input 	ram_block3a35;
input 	ram_block3a3;
input 	ram_block3a36;
input 	ram_block3a4;
input 	ram_block3a37;
input 	ram_block3a5;
input 	ram_block3a38;
input 	ram_block3a6;
input 	ram_block3a39;
input 	ram_block3a7;
input 	ram_block3a40;
input 	ram_block3a8;
input 	ram_block3a41;
input 	ram_block3a9;
input 	ram_block3a42;
input 	ram_block3a10;
input 	ram_block3a43;
input 	ram_block3a11;
input 	ram_block3a44;
input 	ram_block3a12;
input 	ram_block3a45;
input 	ram_block3a13;
input 	ram_block3a46;
input 	ram_block3a14;
input 	ram_block3a47;
input 	ram_block3a15;
input 	ram_block3a48;
input 	ram_block3a16;
input 	ram_block3a49;
input 	ram_block3a17;
input 	ram_block3a50;
input 	ram_block3a18;
input 	ram_block3a51;
input 	ram_block3a19;
input 	ram_block3a52;
input 	ram_block3a20;
input 	ram_block3a53;
input 	ram_block3a21;
input 	ram_block3a54;
input 	ram_block3a22;
input 	ram_block3a55;
input 	ram_block3a23;
input 	ram_block3a56;
input 	ram_block3a24;
input 	ram_block3a57;
input 	ram_block3a25;
input 	ram_block3a58;
input 	ram_block3a26;
input 	ram_block3a59;
input 	ram_block3a27;
input 	ram_block3a60;
input 	ram_block3a28;
input 	ram_block3a61;
input 	ram_block3a29;
input 	ram_block3a62;
input 	ram_block3a30;
input 	ram_block3a63;
input 	ram_block3a31;
output 	is_in_use_reg1;
output 	ram_rom_data_reg_0;
output 	ram_rom_addr_reg_13;
output 	ram_rom_addr_reg_0;
output 	ram_rom_addr_reg_1;
output 	ram_rom_addr_reg_2;
output 	ram_rom_addr_reg_3;
output 	ram_rom_addr_reg_4;
output 	ram_rom_addr_reg_5;
output 	ram_rom_addr_reg_6;
output 	ram_rom_addr_reg_7;
output 	ram_rom_addr_reg_8;
output 	ram_rom_addr_reg_9;
output 	ram_rom_addr_reg_10;
output 	ram_rom_addr_reg_11;
output 	ram_rom_addr_reg_12;
output 	ram_rom_data_reg_1;
output 	ram_rom_data_reg_2;
output 	ram_rom_data_reg_3;
output 	ram_rom_data_reg_4;
output 	ram_rom_data_reg_5;
output 	ram_rom_data_reg_6;
output 	ram_rom_data_reg_7;
output 	ram_rom_data_reg_8;
output 	ram_rom_data_reg_9;
output 	ram_rom_data_reg_10;
output 	ram_rom_data_reg_11;
output 	ram_rom_data_reg_12;
output 	ram_rom_data_reg_13;
output 	ram_rom_data_reg_14;
output 	ram_rom_data_reg_15;
output 	ram_rom_data_reg_16;
output 	ram_rom_data_reg_17;
output 	ram_rom_data_reg_18;
output 	ram_rom_data_reg_19;
output 	ram_rom_data_reg_20;
output 	ram_rom_data_reg_21;
output 	ram_rom_data_reg_22;
output 	ram_rom_data_reg_23;
output 	ram_rom_data_reg_24;
output 	ram_rom_data_reg_25;
output 	ram_rom_data_reg_26;
output 	ram_rom_data_reg_27;
output 	ram_rom_data_reg_28;
output 	ram_rom_data_reg_29;
output 	ram_rom_data_reg_30;
output 	ram_rom_data_reg_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
output 	sdr;
input 	address_reg_b_0;
input 	altera_internal_jtag;
input 	state_4;
input 	[4:0] ir_in;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	raw_tck;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~0_combout ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \ram_rom_data_shift_cntr_reg[0]~6_combout ;
wire \is_in_use_reg~0_combout ;
wire \ram_rom_data_reg[0]~0_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~4_combout ;
wire \ram_rom_data_shift_cntr_reg[1]~5_combout ;
wire \ram_rom_data_shift_cntr_reg[4]~11_combout ;
wire \Add1~3 ;
wire \Add1~4_combout ;
wire \ram_rom_data_shift_cntr_reg[2]~9_combout ;
wire \Add1~5 ;
wire \Add1~6_combout ;
wire \ram_rom_data_shift_cntr_reg[3]~8_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~12_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~10_combout ;
wire \Add1~7 ;
wire \Add1~8_combout ;
wire \ram_rom_data_shift_cntr_reg[4]~7_combout ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \process_0~2_combout ;
wire \ram_rom_data_reg[22]~32_combout ;
wire \ram_rom_addr_reg[0]~15 ;
wire \ram_rom_addr_reg[1]~17 ;
wire \ram_rom_addr_reg[2]~19 ;
wire \ram_rom_addr_reg[3]~21 ;
wire \ram_rom_addr_reg[4]~23 ;
wire \ram_rom_addr_reg[5]~25 ;
wire \ram_rom_addr_reg[6]~27 ;
wire \ram_rom_addr_reg[7]~29 ;
wire \ram_rom_addr_reg[8]~31 ;
wire \ram_rom_addr_reg[9]~33 ;
wire \ram_rom_addr_reg[10]~35 ;
wire \ram_rom_addr_reg[11]~37 ;
wire \ram_rom_addr_reg[12]~39 ;
wire \ram_rom_addr_reg[13]~40_combout ;
wire \process_0~3_combout ;
wire \ram_rom_addr_reg[4]~42_combout ;
wire \ram_rom_addr_reg[4]~43_combout ;
wire \ram_rom_addr_reg[0]~14_combout ;
wire \ram_rom_addr_reg[1]~16_combout ;
wire \ram_rom_addr_reg[2]~18_combout ;
wire \ram_rom_addr_reg[3]~20_combout ;
wire \ram_rom_addr_reg[4]~22_combout ;
wire \ram_rom_addr_reg[5]~24_combout ;
wire \ram_rom_addr_reg[6]~26_combout ;
wire \ram_rom_addr_reg[7]~28_combout ;
wire \ram_rom_addr_reg[8]~30_combout ;
wire \ram_rom_addr_reg[9]~32_combout ;
wire \ram_rom_addr_reg[10]~34_combout ;
wire \ram_rom_addr_reg[11]~36_combout ;
wire \ram_rom_addr_reg[12]~38_combout ;
wire \ram_rom_data_reg[1]~1_combout ;
wire \ram_rom_data_reg[2]~2_combout ;
wire \ram_rom_data_reg[3]~3_combout ;
wire \ram_rom_data_reg[4]~4_combout ;
wire \ram_rom_data_reg[5]~5_combout ;
wire \ram_rom_data_reg[6]~6_combout ;
wire \ram_rom_data_reg[7]~7_combout ;
wire \ram_rom_data_reg[8]~8_combout ;
wire \ram_rom_data_reg[9]~9_combout ;
wire \ram_rom_data_reg[10]~10_combout ;
wire \ram_rom_data_reg[11]~11_combout ;
wire \ram_rom_data_reg[12]~12_combout ;
wire \ram_rom_data_reg[13]~13_combout ;
wire \ram_rom_data_reg[14]~14_combout ;
wire \ram_rom_data_reg[15]~15_combout ;
wire \ram_rom_data_reg[16]~16_combout ;
wire \ram_rom_data_reg[17]~17_combout ;
wire \ram_rom_data_reg[18]~18_combout ;
wire \ram_rom_data_reg[19]~19_combout ;
wire \ram_rom_data_reg[20]~20_combout ;
wire \ram_rom_data_reg[21]~21_combout ;
wire \ram_rom_data_reg[22]~22_combout ;
wire \ram_rom_data_reg[23]~23_combout ;
wire \ram_rom_data_reg[24]~24_combout ;
wire \ram_rom_data_reg[25]~25_combout ;
wire \ram_rom_data_reg[26]~26_combout ;
wire \ram_rom_data_reg[27]~27_combout ;
wire \ram_rom_data_reg[28]~28_combout ;
wire \ram_rom_data_reg[29]~29_combout ;
wire \ram_rom_data_reg[30]~30_combout ;
wire \ram_rom_data_reg[31]~31_combout ;
wire \ir_loaded_address_reg[0]~feeder_combout ;
wire \process_0~0_combout ;
wire \process_0~1_combout ;
wire \ir_loaded_address_reg[1]~feeder_combout ;
wire \ir_loaded_address_reg[2]~feeder_combout ;
wire \bypass_reg_out~0_combout ;
wire \bypass_reg_out~q ;
wire \tdo~0_combout ;
wire [5:0] ram_rom_data_shift_cntr_reg;
wire [3:0] \ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR ;


sld_rom_sr \ram_rom_logic_gen:name_gen:info_rom_sr (
	.WORD_SR_0(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.sdr(sdr),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.TCK(raw_tck),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X43_Y39_N12
cycloneive_lcell_comb \Add1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h55AA;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N20
cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'hC30C;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N22
cycloneive_lcell_comb \Add1~10 (
	.dataa(ram_rom_data_shift_cntr_reg[5]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h5A5A;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X43_Y39_N11
dffeas \ram_rom_data_shift_cntr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[0]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N10
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[0]~6 (
	.dataa(\Add1~0_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[4]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0]~6 .lut_mask = 16'hC0EA;
defparam \ram_rom_data_shift_cntr_reg[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y39_N1
dffeas is_in_use_reg(
	.clk(raw_tck),
	.d(\is_in_use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(ir_in[0]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(is_in_use_reg1),
	.prn(vcc));
// synopsys translate_off
defparam is_in_use_reg.is_wysiwyg = "true";
defparam is_in_use_reg.power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y38_N1
dffeas \ram_rom_data_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[0]~0_combout ),
	.asdata(ram_rom_data_reg_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N27
dffeas \ram_rom_addr_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[13]~40_combout ),
	.asdata(altera_internal_jtag),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N1
dffeas \ram_rom_addr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[0]~14_combout ),
	.asdata(ram_rom_addr_reg_1),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N3
dffeas \ram_rom_addr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[1]~16_combout ),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N5
dffeas \ram_rom_addr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[2]~18_combout ),
	.asdata(ram_rom_addr_reg_3),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N7
dffeas \ram_rom_addr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[3]~20_combout ),
	.asdata(ram_rom_addr_reg_4),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N9
dffeas \ram_rom_addr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[4]~22_combout ),
	.asdata(ram_rom_addr_reg_5),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N11
dffeas \ram_rom_addr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[5]~24_combout ),
	.asdata(ram_rom_addr_reg_6),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N13
dffeas \ram_rom_addr_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[6]~26_combout ),
	.asdata(ram_rom_addr_reg_7),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N15
dffeas \ram_rom_addr_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[7]~28_combout ),
	.asdata(ram_rom_addr_reg_8),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N17
dffeas \ram_rom_addr_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[8]~30_combout ),
	.asdata(ram_rom_addr_reg_9),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N19
dffeas \ram_rom_addr_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[9]~32_combout ),
	.asdata(ram_rom_addr_reg_10),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N21
dffeas \ram_rom_addr_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[10]~34_combout ),
	.asdata(ram_rom_addr_reg_11),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N23
dffeas \ram_rom_addr_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[11]~36_combout ),
	.asdata(ram_rom_addr_reg_12),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N25
dffeas \ram_rom_addr_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[12]~38_combout ),
	.asdata(ram_rom_addr_reg_13),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[4]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y38_N15
dffeas \ram_rom_data_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[1]~1_combout ),
	.asdata(ram_rom_data_reg_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y38_N9
dffeas \ram_rom_data_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[2]~2_combout ),
	.asdata(ram_rom_data_reg_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y38_N31
dffeas \ram_rom_data_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[3]~3_combout ),
	.asdata(ram_rom_data_reg_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y38_N29
dffeas \ram_rom_data_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[4]~4_combout ),
	.asdata(ram_rom_data_reg_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y38_N11
dffeas \ram_rom_data_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[5]~5_combout ),
	.asdata(ram_rom_data_reg_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y38_N5
dffeas \ram_rom_data_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[6]~6_combout ),
	.asdata(ram_rom_data_reg_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X77_Y39_N25
dffeas \ram_rom_data_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[7]~7_combout ),
	.asdata(ram_rom_data_reg_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X77_Y39_N19
dffeas \ram_rom_data_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[8]~8_combout ),
	.asdata(ram_rom_data_reg_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X77_Y39_N9
dffeas \ram_rom_data_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[9]~9_combout ),
	.asdata(ram_rom_data_reg_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X77_Y39_N31
dffeas \ram_rom_data_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[10]~10_combout ),
	.asdata(ram_rom_data_reg_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X77_Y39_N17
dffeas \ram_rom_data_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[11]~11_combout ),
	.asdata(ram_rom_data_reg_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X77_Y39_N23
dffeas \ram_rom_data_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[12]~12_combout ),
	.asdata(ram_rom_data_reg_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X77_Y39_N29
dffeas \ram_rom_data_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[13]~13_combout ),
	.asdata(ram_rom_data_reg_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X77_Y39_N11
dffeas \ram_rom_data_reg[14] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[14]~14_combout ),
	.asdata(ram_rom_data_reg_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_14),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[14] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X77_Y39_N13
dffeas \ram_rom_data_reg[15] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[15]~15_combout ),
	.asdata(ram_rom_data_reg_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_15),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[15] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X77_Y39_N27
dffeas \ram_rom_data_reg[16] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[16]~16_combout ),
	.asdata(ram_rom_data_reg_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_16),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[16] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y43_N9
dffeas \ram_rom_data_reg[17] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[17]~17_combout ),
	.asdata(ram_rom_data_reg_18),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_17),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[17] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y46_N5
dffeas \ram_rom_data_reg[18] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[18]~18_combout ),
	.asdata(ram_rom_data_reg_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_18),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[18] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N13
dffeas \ram_rom_data_reg[19] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[19]~19_combout ),
	.asdata(ram_rom_data_reg_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_19),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[19] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N15
dffeas \ram_rom_data_reg[20] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[20]~20_combout ),
	.asdata(ram_rom_data_reg_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_20),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[20] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N1
dffeas \ram_rom_data_reg[21] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[21]~21_combout ),
	.asdata(ram_rom_data_reg_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_21),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[21] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N27
dffeas \ram_rom_data_reg[22] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[22]~22_combout ),
	.asdata(ram_rom_data_reg_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_22),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[22] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N9
dffeas \ram_rom_data_reg[23] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[23]~23_combout ),
	.asdata(ram_rom_data_reg_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_23),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[23] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N7
dffeas \ram_rom_data_reg[24] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[24]~24_combout ),
	.asdata(ram_rom_data_reg_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_24),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[24] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N17
dffeas \ram_rom_data_reg[25] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[25]~25_combout ),
	.asdata(ram_rom_data_reg_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_25),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[25] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N31
dffeas \ram_rom_data_reg[26] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[26]~26_combout ),
	.asdata(ram_rom_data_reg_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_26),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[26] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N5
dffeas \ram_rom_data_reg[27] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[27]~27_combout ),
	.asdata(ram_rom_data_reg_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_27),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[27] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N11
dffeas \ram_rom_data_reg[28] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[28]~28_combout ),
	.asdata(ram_rom_data_reg_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_28),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[28] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N25
dffeas \ram_rom_data_reg[29] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[29]~29_combout ),
	.asdata(ram_rom_data_reg_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_29),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[29] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y38_N3
dffeas \ram_rom_data_reg[30] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[30]~30_combout ),
	.asdata(ram_rom_data_reg_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_30),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[30] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y38_N5
dffeas \ram_rom_data_reg[31] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[31]~31_combout ),
	.asdata(altera_internal_jtag),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[22]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_31),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[31] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y41_N13
dffeas \ir_loaded_address_reg[0] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[0] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y41_N11
dffeas \ir_loaded_address_reg[1] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[1] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y41_N5
dffeas \ir_loaded_address_reg[2] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[2] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y41_N23
dffeas \ir_loaded_address_reg[3] (
	.clk(raw_tck),
	.d(gnd),
	.asdata(ram_rom_addr_reg_3),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[3] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N22
cycloneive_lcell_comb \tdo~1 (
	.dataa(\tdo~0_combout ),
	.datab(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.datac(gnd),
	.datad(ir_in[0]),
	.cin(gnd),
	.combout(tdo),
	.cout());
// synopsys translate_off
defparam \tdo~1 .lut_mask = 16'hCCAA;
defparam \tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N24
cycloneive_lcell_comb \sdr~0 (
	.dataa(gnd),
	.datab(virtual_ir_scan_reg),
	.datac(node_ena_1),
	.datad(gnd),
	.cin(gnd),
	.combout(sdr),
	.cout());
// synopsys translate_off
defparam \sdr~0 .lut_mask = 16'h3030;
defparam \sdr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N0
cycloneive_lcell_comb \is_in_use_reg~0 (
	.dataa(irf_reg_4_1),
	.datab(gnd),
	.datac(is_in_use_reg1),
	.datad(gnd),
	.cin(gnd),
	.combout(\is_in_use_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \is_in_use_reg~0 .lut_mask = 16'h5050;
defparam \is_in_use_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y38_N0
cycloneive_lcell_comb \ram_rom_data_reg[0]~0 (
	.dataa(ram_block3a0),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a32),
	.cin(gnd),
	.combout(\ram_rom_data_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[0]~0 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N14
cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h3C3F;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N6
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~4 (
	.dataa(irf_reg_1_1),
	.datab(sdr),
	.datac(irf_reg_2_1),
	.datad(state_4),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~4 .lut_mask = 16'hC800;
defparam \ram_rom_data_shift_cntr_reg[5]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N8
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[1]~5 (
	.dataa(\Equal1~1_combout ),
	.datab(\Add1~2_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1]~5 .lut_mask = 16'h4C50;
defparam \ram_rom_data_shift_cntr_reg[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N9
dffeas \ram_rom_data_shift_cntr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[1]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N4
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[4]~11 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(\Equal1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[4]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4]~11 .lut_mask = 16'h007F;
defparam \ram_rom_data_shift_cntr_reg[4]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N16
cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'hC30C;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N28
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[2]~9 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[4]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[2]),
	.datad(\Add1~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2]~9 .lut_mask = 16'hD5C0;
defparam \ram_rom_data_shift_cntr_reg[2]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N29
dffeas \ram_rom_data_shift_cntr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[2]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N18
cycloneive_lcell_comb \Add1~6 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h3C3F;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N2
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[3]~8 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[4]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[3]),
	.datad(\Add1~6_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3]~8 .lut_mask = 16'hD5C0;
defparam \ram_rom_data_shift_cntr_reg[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N3
dffeas \ram_rom_data_shift_cntr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[3]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N6
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~12 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(\Equal1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~12 .lut_mask = 16'h80FF;
defparam \ram_rom_data_shift_cntr_reg[5]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N26
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~10 (
	.dataa(\Add1~10_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[4]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~10 .lut_mask = 16'hC0EA;
defparam \ram_rom_data_shift_cntr_reg[5]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N27
dffeas \ram_rom_data_shift_cntr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[5]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N0
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[4]~7 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[4]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[4]),
	.datad(\Add1~8_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4]~7 .lut_mask = 16'hD5C0;
defparam \ram_rom_data_shift_cntr_reg[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N1
dffeas \ram_rom_data_shift_cntr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[4]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N24
cycloneive_lcell_comb \Equal1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[2]),
	.datab(ram_rom_data_shift_cntr_reg[3]),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(ram_rom_data_shift_cntr_reg[4]),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h0800;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N30
cycloneive_lcell_comb \Equal1~1 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'hAA00;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N8
cycloneive_lcell_comb \process_0~2 (
	.dataa(\Equal1~1_combout ),
	.datab(ir_in[3]),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\process_0~2_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~2 .lut_mask = 16'h1333;
defparam \process_0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N16
cycloneive_lcell_comb \ram_rom_data_reg[22]~32 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\process_0~2_combout ),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_reg[22]~32_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[22]~32 .lut_mask = 16'hFF0F;
defparam \ram_rom_data_reg[22]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N0
cycloneive_lcell_comb \ram_rom_addr_reg[0]~14 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[0]~14_combout ),
	.cout(\ram_rom_addr_reg[0]~15 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[0]~14 .lut_mask = 16'h33CC;
defparam \ram_rom_addr_reg[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N2
cycloneive_lcell_comb \ram_rom_addr_reg[1]~16 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[0]~15 ),
	.combout(\ram_rom_addr_reg[1]~16_combout ),
	.cout(\ram_rom_addr_reg[1]~17 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[1]~16 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[1]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N4
cycloneive_lcell_comb \ram_rom_addr_reg[2]~18 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[1]~17 ),
	.combout(\ram_rom_addr_reg[2]~18_combout ),
	.cout(\ram_rom_addr_reg[2]~19 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[2]~18 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[2]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N6
cycloneive_lcell_comb \ram_rom_addr_reg[3]~20 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[2]~19 ),
	.combout(\ram_rom_addr_reg[3]~20_combout ),
	.cout(\ram_rom_addr_reg[3]~21 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[3]~20 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[3]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N8
cycloneive_lcell_comb \ram_rom_addr_reg[4]~22 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[3]~21 ),
	.combout(\ram_rom_addr_reg[4]~22_combout ),
	.cout(\ram_rom_addr_reg[4]~23 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[4]~22 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[4]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N10
cycloneive_lcell_comb \ram_rom_addr_reg[5]~24 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[4]~23 ),
	.combout(\ram_rom_addr_reg[5]~24_combout ),
	.cout(\ram_rom_addr_reg[5]~25 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~24 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[5]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N12
cycloneive_lcell_comb \ram_rom_addr_reg[6]~26 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[5]~25 ),
	.combout(\ram_rom_addr_reg[6]~26_combout ),
	.cout(\ram_rom_addr_reg[6]~27 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[6]~26 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[6]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N14
cycloneive_lcell_comb \ram_rom_addr_reg[7]~28 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[6]~27 ),
	.combout(\ram_rom_addr_reg[7]~28_combout ),
	.cout(\ram_rom_addr_reg[7]~29 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[7]~28 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[7]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N16
cycloneive_lcell_comb \ram_rom_addr_reg[8]~30 (
	.dataa(ram_rom_addr_reg_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[7]~29 ),
	.combout(\ram_rom_addr_reg[8]~30_combout ),
	.cout(\ram_rom_addr_reg[8]~31 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[8]~30 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[8]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N18
cycloneive_lcell_comb \ram_rom_addr_reg[9]~32 (
	.dataa(ram_rom_addr_reg_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[8]~31 ),
	.combout(\ram_rom_addr_reg[9]~32_combout ),
	.cout(\ram_rom_addr_reg[9]~33 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[9]~32 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[9]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N20
cycloneive_lcell_comb \ram_rom_addr_reg[10]~34 (
	.dataa(ram_rom_addr_reg_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[9]~33 ),
	.combout(\ram_rom_addr_reg[10]~34_combout ),
	.cout(\ram_rom_addr_reg[10]~35 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[10]~34 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[10]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N22
cycloneive_lcell_comb \ram_rom_addr_reg[11]~36 (
	.dataa(ram_rom_addr_reg_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[10]~35 ),
	.combout(\ram_rom_addr_reg[11]~36_combout ),
	.cout(\ram_rom_addr_reg[11]~37 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[11]~36 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[11]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N24
cycloneive_lcell_comb \ram_rom_addr_reg[12]~38 (
	.dataa(ram_rom_addr_reg_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[11]~37 ),
	.combout(\ram_rom_addr_reg[12]~38_combout ),
	.cout(\ram_rom_addr_reg[12]~39 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[12]~38 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[12]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N26
cycloneive_lcell_comb \ram_rom_addr_reg[13]~40 (
	.dataa(ram_rom_addr_reg_13),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\ram_rom_addr_reg[12]~39 ),
	.combout(\ram_rom_addr_reg[13]~40_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[13]~40 .lut_mask = 16'h5A5A;
defparam \ram_rom_addr_reg[13]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N30
cycloneive_lcell_comb \process_0~3 (
	.dataa(node_ena_1),
	.datab(ir_in[3]),
	.datac(virtual_ir_scan_reg),
	.datad(state_4),
	.cin(gnd),
	.combout(\process_0~3_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~3 .lut_mask = 16'h0800;
defparam \process_0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N4
cycloneive_lcell_comb \ram_rom_addr_reg[4]~42 (
	.dataa(\Equal1~1_combout ),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(\process_0~3_combout ),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[4]~42_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[4]~42 .lut_mask = 16'hF2F0;
defparam \ram_rom_addr_reg[4]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N18
cycloneive_lcell_comb \ram_rom_addr_reg[4]~43 (
	.dataa(irf_reg_2_1),
	.datab(state_8),
	.datac(\ram_rom_addr_reg[4]~42_combout ),
	.datad(sdr),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[4]~43_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[4]~43 .lut_mask = 16'hF8F0;
defparam \ram_rom_addr_reg[4]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y38_N14
cycloneive_lcell_comb \ram_rom_data_reg[1]~1 (
	.dataa(ram_block3a33),
	.datab(ram_block3a1),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[1]~1 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y38_N8
cycloneive_lcell_comb \ram_rom_data_reg[2]~2 (
	.dataa(ram_block3a2),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a34),
	.cin(gnd),
	.combout(\ram_rom_data_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[2]~2 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y38_N30
cycloneive_lcell_comb \ram_rom_data_reg[3]~3 (
	.dataa(ram_block3a3),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a35),
	.cin(gnd),
	.combout(\ram_rom_data_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[3]~3 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y38_N28
cycloneive_lcell_comb \ram_rom_data_reg[4]~4 (
	.dataa(ram_block3a36),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a4),
	.cin(gnd),
	.combout(\ram_rom_data_reg[4]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[4]~4 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y38_N10
cycloneive_lcell_comb \ram_rom_data_reg[5]~5 (
	.dataa(ram_block3a5),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a37),
	.cin(gnd),
	.combout(\ram_rom_data_reg[5]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[5]~5 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y38_N4
cycloneive_lcell_comb \ram_rom_data_reg[6]~6 (
	.dataa(ram_block3a38),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a6),
	.cin(gnd),
	.combout(\ram_rom_data_reg[6]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[6]~6 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y39_N24
cycloneive_lcell_comb \ram_rom_data_reg[7]~7 (
	.dataa(ram_block3a7),
	.datab(ram_block3a39),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[7]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[7]~7 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y39_N18
cycloneive_lcell_comb \ram_rom_data_reg[8]~8 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a40),
	.datac(gnd),
	.datad(ram_block3a8),
	.cin(gnd),
	.combout(\ram_rom_data_reg[8]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[8]~8 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y39_N8
cycloneive_lcell_comb \ram_rom_data_reg[9]~9 (
	.dataa(ram_block3a9),
	.datab(ram_block3a41),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[9]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[9]~9 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y39_N30
cycloneive_lcell_comb \ram_rom_data_reg[10]~10 (
	.dataa(ram_block3a42),
	.datab(ram_block3a10),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[10]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[10]~10 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y39_N16
cycloneive_lcell_comb \ram_rom_data_reg[11]~11 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a11),
	.datac(gnd),
	.datad(ram_block3a43),
	.cin(gnd),
	.combout(\ram_rom_data_reg[11]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[11]~11 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y39_N22
cycloneive_lcell_comb \ram_rom_data_reg[12]~12 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a12),
	.datac(gnd),
	.datad(ram_block3a44),
	.cin(gnd),
	.combout(\ram_rom_data_reg[12]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[12]~12 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y39_N28
cycloneive_lcell_comb \ram_rom_data_reg[13]~13 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a45),
	.datac(gnd),
	.datad(ram_block3a13),
	.cin(gnd),
	.combout(\ram_rom_data_reg[13]~13_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[13]~13 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y39_N10
cycloneive_lcell_comb \ram_rom_data_reg[14]~14 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a46),
	.datac(gnd),
	.datad(ram_block3a14),
	.cin(gnd),
	.combout(\ram_rom_data_reg[14]~14_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[14]~14 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y39_N12
cycloneive_lcell_comb \ram_rom_data_reg[15]~15 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a15),
	.datac(gnd),
	.datad(ram_block3a47),
	.cin(gnd),
	.combout(\ram_rom_data_reg[15]~15_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[15]~15 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y39_N26
cycloneive_lcell_comb \ram_rom_data_reg[16]~16 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a16),
	.datac(gnd),
	.datad(ram_block3a48),
	.cin(gnd),
	.combout(\ram_rom_data_reg[16]~16_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[16]~16 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y43_N8
cycloneive_lcell_comb \ram_rom_data_reg[17]~17 (
	.dataa(ram_block3a49),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a17),
	.cin(gnd),
	.combout(\ram_rom_data_reg[17]~17_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[17]~17 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y46_N4
cycloneive_lcell_comb \ram_rom_data_reg[18]~18 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a50),
	.datac(gnd),
	.datad(ram_block3a18),
	.cin(gnd),
	.combout(\ram_rom_data_reg[18]~18_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[18]~18 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N12
cycloneive_lcell_comb \ram_rom_data_reg[19]~19 (
	.dataa(ram_block3a51),
	.datab(ram_block3a19),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[19]~19_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[19]~19 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N14
cycloneive_lcell_comb \ram_rom_data_reg[20]~20 (
	.dataa(ram_block3a52),
	.datab(ram_block3a20),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[20]~20_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[20]~20 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N0
cycloneive_lcell_comb \ram_rom_data_reg[21]~21 (
	.dataa(ram_block3a53),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a21),
	.cin(gnd),
	.combout(\ram_rom_data_reg[21]~21_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[21]~21 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N26
cycloneive_lcell_comb \ram_rom_data_reg[22]~22 (
	.dataa(ram_block3a22),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a54),
	.cin(gnd),
	.combout(\ram_rom_data_reg[22]~22_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[22]~22 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N8
cycloneive_lcell_comb \ram_rom_data_reg[23]~23 (
	.dataa(ram_block3a55),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a23),
	.cin(gnd),
	.combout(\ram_rom_data_reg[23]~23_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[23]~23 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N6
cycloneive_lcell_comb \ram_rom_data_reg[24]~24 (
	.dataa(ram_block3a56),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a24),
	.cin(gnd),
	.combout(\ram_rom_data_reg[24]~24_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[24]~24 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N16
cycloneive_lcell_comb \ram_rom_data_reg[25]~25 (
	.dataa(ram_block3a25),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a57),
	.cin(gnd),
	.combout(\ram_rom_data_reg[25]~25_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[25]~25 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N30
cycloneive_lcell_comb \ram_rom_data_reg[26]~26 (
	.dataa(ram_block3a26),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a58),
	.cin(gnd),
	.combout(\ram_rom_data_reg[26]~26_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[26]~26 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N4
cycloneive_lcell_comb \ram_rom_data_reg[27]~27 (
	.dataa(ram_block3a59),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a27),
	.cin(gnd),
	.combout(\ram_rom_data_reg[27]~27_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[27]~27 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N10
cycloneive_lcell_comb \ram_rom_data_reg[28]~28 (
	.dataa(ram_block3a28),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a60),
	.cin(gnd),
	.combout(\ram_rom_data_reg[28]~28_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[28]~28 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N24
cycloneive_lcell_comb \ram_rom_data_reg[29]~29 (
	.dataa(ram_block3a61),
	.datab(ram_block3a29),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[29]~29_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[29]~29 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y38_N2
cycloneive_lcell_comb \ram_rom_data_reg[30]~30 (
	.dataa(ram_block3a30),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a62),
	.cin(gnd),
	.combout(\ram_rom_data_reg[30]~30_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[30]~30 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N4
cycloneive_lcell_comb \ram_rom_data_reg[31]~31 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a31),
	.datac(gnd),
	.datad(ram_block3a63),
	.cin(gnd),
	.combout(\ram_rom_data_reg[31]~31_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[31]~31 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y41_N12
cycloneive_lcell_comb \ir_loaded_address_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_0),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y41_N24
cycloneive_lcell_comb \process_0~0 (
	.dataa(gnd),
	.datab(irf_reg_4_1),
	.datac(ir_in[0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\process_0~0_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~0 .lut_mask = 16'hFCFC;
defparam \process_0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N26
cycloneive_lcell_comb \process_0~1 (
	.dataa(node_ena_1),
	.datab(virtual_ir_scan_reg),
	.datac(state_5),
	.datad(ir_in[3]),
	.cin(gnd),
	.combout(\process_0~1_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~1 .lut_mask = 16'h2000;
defparam \process_0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y41_N10
cycloneive_lcell_comb \ir_loaded_address_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_1),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y41_N4
cycloneive_lcell_comb \ir_loaded_address_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_2),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N10
cycloneive_lcell_comb \bypass_reg_out~0 (
	.dataa(node_ena_1),
	.datab(altera_internal_jtag),
	.datac(\bypass_reg_out~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\bypass_reg_out~0_combout ),
	.cout());
// synopsys translate_off
defparam \bypass_reg_out~0 .lut_mask = 16'hD8D8;
defparam \bypass_reg_out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y39_N11
dffeas bypass_reg_out(
	.clk(raw_tck),
	.d(\bypass_reg_out~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\bypass_reg_out~q ),
	.prn(vcc));
// synopsys translate_off
defparam bypass_reg_out.is_wysiwyg = "true";
defparam bypass_reg_out.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y39_N12
cycloneive_lcell_comb \tdo~0 (
	.dataa(\bypass_reg_out~q ),
	.datab(ram_rom_data_reg_0),
	.datac(irf_reg_2_1),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \tdo~0 .lut_mask = 16'hCCCA;
defparam \tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_rom_sr (
	WORD_SR_0,
	sdr,
	altera_internal_jtag,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	TCK,
	devpor,
	devclrn,
	devoe);
output 	WORD_SR_0;
input 	sdr;
input 	altera_internal_jtag;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	TCK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \WORD_SR~3_combout ;
wire \WORD_SR~7_combout ;
wire \WORD_SR~8_combout ;
wire \WORD_SR~10_combout ;
wire \WORD_SR~11_combout ;
wire \WORD_SR~13_combout ;
wire \WORD_SR~14_combout ;
wire \clear_signal~combout ;
wire \WORD_SR~15_combout ;
wire \WORD_SR[2]~6_combout ;
wire \WORD_SR~12_combout ;
wire \WORD_SR~9_combout ;
wire \word_counter[0]~7_combout ;
wire \word_counter[3]~15_combout ;
wire \word_counter[4]~14_combout ;
wire \word_counter[4]~13_combout ;
wire \word_counter[4]~19_combout ;
wire \word_counter[0]~8 ;
wire \word_counter[1]~9_combout ;
wire \word_counter[1]~10 ;
wire \word_counter[2]~11_combout ;
wire \word_counter[2]~12 ;
wire \word_counter[3]~16 ;
wire \word_counter[4]~17_combout ;
wire \WORD_SR~2_combout ;
wire \WORD_SR~4_combout ;
wire \WORD_SR~5_combout ;
wire [4:0] word_counter;
wire [3:0] WORD_SR;


// Location: LCCOMB_X41_Y39_N10
cycloneive_lcell_comb \WORD_SR~3 (
	.dataa(word_counter[0]),
	.datab(word_counter[4]),
	.datac(word_counter[1]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\WORD_SR~3_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~3 .lut_mask = 16'hD0C4;
defparam \WORD_SR~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N8
cycloneive_lcell_comb \WORD_SR~7 (
	.dataa(word_counter[0]),
	.datab(word_counter[1]),
	.datac(word_counter[4]),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~7 .lut_mask = 16'h0045;
defparam \WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N10
cycloneive_lcell_comb \WORD_SR~8 (
	.dataa(gnd),
	.datab(word_counter[3]),
	.datac(\WORD_SR~7_combout ),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~8 .lut_mask = 16'h0030;
defparam \WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y39_N2
cycloneive_lcell_comb \WORD_SR~10 (
	.dataa(word_counter[0]),
	.datab(word_counter[4]),
	.datac(word_counter[1]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~10 .lut_mask = 16'hADCC;
defparam \WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y39_N12
cycloneive_lcell_comb \WORD_SR~11 (
	.dataa(gnd),
	.datab(\WORD_SR~10_combout ),
	.datac(\WORD_SR~2_combout ),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~11 .lut_mask = 16'hCC30;
defparam \WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N28
cycloneive_lcell_comb \WORD_SR~13 (
	.dataa(word_counter[1]),
	.datab(word_counter[3]),
	.datac(word_counter[4]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~13 .lut_mask = 16'h0800;
defparam \WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N26
cycloneive_lcell_comb \WORD_SR~14 (
	.dataa(word_counter[0]),
	.datab(\WORD_SR~13_combout ),
	.datac(altera_internal_jtag),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~14 .lut_mask = 16'hF044;
defparam \WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y39_N25
dffeas \WORD_SR[0] (
	.clk(TCK),
	.d(\WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR_0),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[0] .is_wysiwyg = "true";
defparam \WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N20
cycloneive_lcell_comb clear_signal(
	.dataa(gnd),
	.datab(gnd),
	.datac(state_8),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam clear_signal.lut_mask = 16'hF000;
defparam clear_signal.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N22
cycloneive_lcell_comb \WORD_SR~15 (
	.dataa(\WORD_SR~14_combout ),
	.datab(gnd),
	.datac(state_8),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\WORD_SR~15_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~15 .lut_mask = 16'h0AAA;
defparam \WORD_SR~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N2
cycloneive_lcell_comb \WORD_SR[2]~6 (
	.dataa(state_3),
	.datab(\clear_signal~combout ),
	.datac(sdr),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR[2]~6_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR[2]~6 .lut_mask = 16'hFCEC;
defparam \WORD_SR[2]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y39_N23
dffeas \WORD_SR[3] (
	.clk(TCK),
	.d(\WORD_SR~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[3]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[3] .is_wysiwyg = "true";
defparam \WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N4
cycloneive_lcell_comb \WORD_SR~12 (
	.dataa(\WORD_SR~11_combout ),
	.datab(\clear_signal~combout ),
	.datac(WORD_SR[3]),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~12 .lut_mask = 16'h3022;
defparam \WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y39_N5
dffeas \WORD_SR[2] (
	.clk(TCK),
	.d(\WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[2]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[2] .is_wysiwyg = "true";
defparam \WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N6
cycloneive_lcell_comb \WORD_SR~9 (
	.dataa(\WORD_SR~8_combout ),
	.datab(\clear_signal~combout ),
	.datac(WORD_SR[2]),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~9 .lut_mask = 16'h3222;
defparam \WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y39_N7
dffeas \WORD_SR[1] (
	.clk(TCK),
	.d(\WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[2]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[1]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[1] .is_wysiwyg = "true";
defparam \WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y39_N16
cycloneive_lcell_comb \word_counter[0]~7 (
	.dataa(gnd),
	.datab(word_counter[0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\word_counter[0]~7_combout ),
	.cout(\word_counter[0]~8 ));
// synopsys translate_off
defparam \word_counter[0]~7 .lut_mask = 16'h33CC;
defparam \word_counter[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y39_N22
cycloneive_lcell_comb \word_counter[3]~15 (
	.dataa(word_counter[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[2]~12 ),
	.combout(\word_counter[3]~15_combout ),
	.cout(\word_counter[3]~16 ));
// synopsys translate_off
defparam \word_counter[3]~15 .lut_mask = 16'h5A5F;
defparam \word_counter[3]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N12
cycloneive_lcell_comb \word_counter[4]~14 (
	.dataa(state_3),
	.datab(\clear_signal~combout ),
	.datac(sdr),
	.datad(state_4),
	.cin(gnd),
	.combout(\word_counter[4]~14_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~14 .lut_mask = 16'hCCEC;
defparam \word_counter[4]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y39_N23
dffeas \word_counter[3] (
	.clk(TCK),
	.d(\word_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[4]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[4]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[3]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[3] .is_wysiwyg = "true";
defparam \word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N18
cycloneive_lcell_comb \word_counter[4]~13 (
	.dataa(word_counter[1]),
	.datab(word_counter[3]),
	.datac(word_counter[4]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\word_counter[4]~13_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~13 .lut_mask = 16'hEFFF;
defparam \word_counter[4]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N0
cycloneive_lcell_comb \word_counter[4]~19 (
	.dataa(state_8),
	.datab(\word_counter[4]~13_combout ),
	.datac(word_counter[0]),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\word_counter[4]~19_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~19 .lut_mask = 16'hAB03;
defparam \word_counter[4]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y39_N17
dffeas \word_counter[0] (
	.clk(TCK),
	.d(\word_counter[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[4]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[4]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[0]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[0] .is_wysiwyg = "true";
defparam \word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y39_N18
cycloneive_lcell_comb \word_counter[1]~9 (
	.dataa(gnd),
	.datab(word_counter[1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[0]~8 ),
	.combout(\word_counter[1]~9_combout ),
	.cout(\word_counter[1]~10 ));
// synopsys translate_off
defparam \word_counter[1]~9 .lut_mask = 16'h3C3F;
defparam \word_counter[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X41_Y39_N19
dffeas \word_counter[1] (
	.clk(TCK),
	.d(\word_counter[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[4]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[4]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[1]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[1] .is_wysiwyg = "true";
defparam \word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y39_N20
cycloneive_lcell_comb \word_counter[2]~11 (
	.dataa(gnd),
	.datab(word_counter[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[1]~10 ),
	.combout(\word_counter[2]~11_combout ),
	.cout(\word_counter[2]~12 ));
// synopsys translate_off
defparam \word_counter[2]~11 .lut_mask = 16'hC30C;
defparam \word_counter[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X41_Y39_N21
dffeas \word_counter[2] (
	.clk(TCK),
	.d(\word_counter[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[4]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[4]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[2]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[2] .is_wysiwyg = "true";
defparam \word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y39_N24
cycloneive_lcell_comb \word_counter[4]~17 (
	.dataa(gnd),
	.datab(word_counter[4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\word_counter[3]~16 ),
	.combout(\word_counter[4]~17_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~17 .lut_mask = 16'hC3C3;
defparam \word_counter[4]~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X41_Y39_N25
dffeas \word_counter[4] (
	.clk(TCK),
	.d(\word_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[4]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[4]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[4]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[4] .is_wysiwyg = "true";
defparam \word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y39_N8
cycloneive_lcell_comb \WORD_SR~2 (
	.dataa(word_counter[1]),
	.datab(word_counter[4]),
	.datac(word_counter[3]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\WORD_SR~2_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~2 .lut_mask = 16'h3005;
defparam \WORD_SR~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y39_N0
cycloneive_lcell_comb \WORD_SR~4 (
	.dataa(\WORD_SR~3_combout ),
	.datab(gnd),
	.datac(\WORD_SR~2_combout ),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~4_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~4 .lut_mask = 16'hAAA0;
defparam \WORD_SR~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N24
cycloneive_lcell_comb \WORD_SR~5 (
	.dataa(WORD_SR[1]),
	.datab(\clear_signal~combout ),
	.datac(\WORD_SR~4_combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~5_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~5 .lut_mask = 16'h2230;
defparam \WORD_SR~5 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule
