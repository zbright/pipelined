`include "datapath_cache_if.vh"
`include "cpu_types_pkg.vh"

module request_unit (
	input logic CLK,
	input logic dhit,
	input logic request_dmemREN,
	input logic request_dmemWEN,
	output logic request_dmemREN_output,
	output logic request_dmemWEN_output	
	);

	import cpu_types_pkg::*;

	//assign request_dmemREN_output = dhit ? 0 : request_dmemREN;
	//assign request_dmemWEN_output = dhit ? 0 : request_dmemWEN;

	
	always_ff@(posedge CLK)
	begin
		//not sure where to put it
		request_dmemREN_output = request_dmemREN;
		request_dmemWEN_output = request_dmemWEN;
		if (dhit == 1) begin
			request_dmemREN_output = 0;
			request_dmemWEN_output = 0;
		end else begin
			request_dmemREN_output = request_dmemREN;
			request_dmemWEN_output = request_dmemWEN;
		end
	end

endmodule
		
