module alu_fpga (
	input logic [3:0] KEY,
	input logic [17:0] SW,
	output logic [17:0] LEDR,
	output logic [6:0]HEX0,
	output logic [6:0]HEX1,
	output logic [6:0]HEX2,
	output logic [6:0]HEX3,
	output logic [6:0]HEX4,
	output logic [6:0]HEX5,
	output logic [6:0]HEX6,
	output logic [6:0]HEX7
);

logic [31:0] TEMPA;
logic [31:0] TEMPB;
logic [31:0] OUTPUT;
logic [14:0] SWITCHVAL;
logic [3:0] OPCODE;
logic ABSELECT;
logic TOGGLE;

assign SWITCHVAL = SW[14:0];
assign ABSELECT = SW[17];
assign TOGGLE = SW[15];
assign OPCODE = KEY[3:0];
assign LEDR[0] = NEGATIVE;
assign LEDR[1] = OVERFLOW;
assign LEDR[2] = ZERO;
//assign LEDR[3] = OPCODE[1];
//assign LEDR[4] = OPCODE[2];
//assign LEDR[5] = OPCODE[3];

//assigning values
assign TEMPA [14:0] = ABSELECT ? SWITCHVAL : TEMPA;
assign TEMPB [14:0] = ABSELECT ? TEMPB : SWITCHVAL;
//filling in values for a
assign TEMPA [15] = TOGGLE ? 1 : 0;
assign TEMPA [16] = TOGGLE ? 1 : 0;
assign TEMPA [17] = TOGGLE ? 1 : 0;
assign TEMPA [18] = TOGGLE ? 1 : 0;
assign TEMPA [19] = TOGGLE ? 1 : 0;
assign TEMPA [20] = TOGGLE ? 1 : 0;
assign TEMPA [21] = TOGGLE ? 1 : 0;
assign TEMPA [22] = TOGGLE ? 1 : 0;
assign TEMPA [23] = TOGGLE ? 1 : 0;
assign TEMPA [24] = TOGGLE ? 1 : 0;
assign TEMPA [25] = TOGGLE ? 1 : 0;
assign TEMPA [26] = TOGGLE ? 1 : 0;
assign TEMPA [27] = TOGGLE ? 1 : 0;
assign TEMPA [28] = TOGGLE ? 1 : 0;
assign TEMPA [29] = TOGGLE ? 1 : 0;
assign TEMPA [30] = TOGGLE ? 1 : 0;
assign TEMPA [31] = TOGGLE ? 1 : 0;
//filling in values for b
assign TEMPB [15] = TOGGLE ? 1 : 0;
assign TEMPB [16] = TOGGLE ? 1 : 0;
assign TEMPB [17] = TOGGLE ? 1 : 0;
assign TEMPB [18] = TOGGLE ? 1 : 0;
assign TEMPB [19] = TOGGLE ? 1 : 0;
assign TEMPB [20] = TOGGLE ? 1 : 0;
assign TEMPB [21] = TOGGLE ? 1 : 0;
assign TEMPB [22] = TOGGLE ? 1 : 0;
assign TEMPB [23] = TOGGLE ? 1 : 0;
assign TEMPB [24] = TOGGLE ? 1 : 0;
assign TEMPB [25] = TOGGLE ? 1 : 0;
assign TEMPB [26] = TOGGLE ? 1 : 0;
assign TEMPB [27] = TOGGLE ? 1 : 0;
assign TEMPB [28] = TOGGLE ? 1 : 0;
assign TEMPB [29] = TOGGLE ? 1 : 0;
assign TEMPB [30] = TOGGLE ? 1 : 0;
assign TEMPB [31] = TOGGLE ? 1 : 0;

  always_comb
  begin
    unique casez (OUTPUT[3:0])
      'h0: HEX0 = 7'b1000000;
      'h1: HEX0 = 7'b1111001;
      'h2: HEX0 = 7'b0100100;
      'h3: HEX0 = 7'b0110000;
      'h4: HEX0 = 7'b0011001;
      'h5: HEX0 = 7'b0010010;
      'h6: HEX0 = 7'b0000010;
      'h7: HEX0 = 7'b1111000;
      'h8: HEX0 = 7'b0000000;
      'h9: HEX0 = 7'b0010000;
      'ha: HEX0 = 7'b0001000;
      'hb: HEX0 = 7'b0000011;
      'hc: HEX0 = 7'b0100111;
      'hd: HEX0 = 7'b0100001;
      'he: HEX0 = 7'b0000110;
      'hf: HEX0 = 7'b0001110;
    endcase
    
    unique casez (OUTPUT[7:4])
      'h0: HEX1 = 7'b1000000;
      'h1: HEX1 = 7'b1111001;
      'h2: HEX1 = 7'b0100100;
      'h3: HEX1 = 7'b0110000;
      'h4: HEX1 = 7'b0011001;
      'h5: HEX1 = 7'b0010010;
      'h6: HEX1 = 7'b0000010;
      'h7: HEX1 = 7'b1111000;
      'h8: HEX1 = 7'b0000000;
      'h9: HEX1 = 7'b0010000;
      'ha: HEX1 = 7'b0001000;
      'hb: HEX1 = 7'b0000011;
      'hc: HEX1 = 7'b0100111;
      'hd: HEX1 = 7'b0100001;
      'he: HEX1 = 7'b0000110;
      'hf: HEX1 = 7'b0001110;
    endcase

    unique casez (OUTPUT[11:8])
      'h0: HEX2 = 7'b1000000;
      'h1: HEX2 = 7'b1111001;
      'h2: HEX2 = 7'b0100100;
      'h3: HEX2 = 7'b0110000;
      'h4: HEX2 = 7'b0011001;
      'h5: HEX2 = 7'b0010010;
      'h6: HEX2 = 7'b0000010;
      'h7: HEX2 = 7'b1111000;
      'h8: HEX2 = 7'b0000000;
      'h9: HEX2 = 7'b0010000;
      'ha: HEX2 = 7'b0001000;
      'hb: HEX2 = 7'b0000011;
      'hc: HEX2 = 7'b0100111;
      'hd: HEX2 = 7'b0100001;
      'he: HEX2 = 7'b0000110;
      'hf: HEX2 = 7'b0001110;
    endcase

    unique casez (OUTPUT[15:12])
      'h0: HEX3 = 7'b1000000;
      'h1: HEX3 = 7'b1111001;
      'h2: HEX3 = 7'b0100100;
      'h3: HEX3 = 7'b0110000;
      'h4: HEX3 = 7'b0011001;
      'h5: HEX3 = 7'b0010010;
      'h6: HEX3 = 7'b0000010;
      'h7: HEX3 = 7'b1111000;
      'h8: HEX3 = 7'b0000000;
      'h9: HEX3 = 7'b0010000;
      'ha: HEX3 = 7'b0001000;
      'hb: HEX3 = 7'b0000011;
      'hc: HEX3 = 7'b0100111;
      'hd: HEX3 = 7'b0100001;
      'he: HEX3 = 7'b0000110;
      'hf: HEX3 = 7'b0001110;
    endcase

    unique casez (OUTPUT[19:16])
      'h0: HEX4 = 7'b1000000;
      'h1: HEX4 = 7'b1111001;
      'h2: HEX4 = 7'b0100100;
      'h3: HEX4 = 7'b0110000;
      'h4: HEX4 = 7'b0011001;
      'h5: HEX4 = 7'b0010010;
      'h6: HEX4 = 7'b0000010;
      'h7: HEX4 = 7'b1111000;
      'h8: HEX4 = 7'b0000000;
      'h9: HEX4 = 7'b0010000;
      'ha: HEX4 = 7'b0001000;
      'hb: HEX4 = 7'b0000011;
      'hc: HEX4 = 7'b0100111;
      'hd: HEX4 = 7'b0100001;
      'he: HEX4 = 7'b0000110;
      'hf: HEX4 = 7'b0001110;
    endcase

    unique casez (OUTPUT[23:20])
      'h0: HEX5 = 7'b1000000;
      'h1: HEX5 = 7'b1111001;
      'h2: HEX5 = 7'b0100100;
      'h3: HEX5 = 7'b0110000;
      'h4: HEX5 = 7'b0011001;
      'h5: HEX5 = 7'b0010010;
      'h6: HEX5 = 7'b0000010;
      'h7: HEX5 = 7'b1111000;
      'h8: HEX5 = 7'b0000000;
      'h9: HEX5 = 7'b0010000;
      'ha: HEX5 = 7'b0001000;
      'hb: HEX5 = 7'b0000011;
      'hc: HEX5 = 7'b0100111;
      'hd: HEX5 = 7'b0100001;
      'he: HEX5 = 7'b0000110;
      'hf: HEX5 = 7'b0001110;
    endcase

    unique casez (OUTPUT[27:24])
      'h0: HEX6 = 7'b1000000;
      'h1: HEX6 = 7'b1111001;
      'h2: HEX6 = 7'b0100100;
      'h3: HEX6 = 7'b0110000;
      'h4: HEX6 = 7'b0011001;
      'h5: HEX6 = 7'b0010010;
      'h6: HEX6 = 7'b0000010;
      'h7: HEX6 = 7'b1111000;
      'h8: HEX6 = 7'b0000000;
      'h9: HEX6 = 7'b0010000;
      'ha: HEX6 = 7'b0001000;
      'hb: HEX6 = 7'b0000011;
      'hc: HEX6 = 7'b0100111;
      'hd: HEX6 = 7'b0100001;
      'he: HEX6 = 7'b0000110;
      'hf: HEX6 = 7'b0001110;
    endcase

    unique casez (OUTPUT[31:28])
      'h0: HEX7 = 7'b1000000;
      'h1: HEX7 = 7'b1111001;
      'h2: HEX7 = 7'b0100100;
      'h3: HEX7 = 7'b0110000;
      'h4: HEX7 = 7'b0011001;
      'h5: HEX7 = 7'b0010010;
      'h6: HEX7 = 7'b0000010;
      'h7: HEX7 = 7'b1111000;
      'h8: HEX7 = 7'b0000000;
      'h9: HEX7 = 7'b0010000;
      'ha: HEX7 = 7'b0001000;
      'hb: HEX7 = 7'b0000011;
      'hc: HEX7 = 7'b0100111;
      'hd: HEX7 = 7'b0100001;
      'he: HEX7 = 7'b0000110;
      'hf: HEX7 = 7'b0001110;
    endcase
	
  end

 alu ALU(TEMPA, TEMPB, OPCODE, OUTPUT, NEGATIVE, OVERFLOW, ZERO);

//just a test

/*assign rfif.wsel = SW[4:0];
assign rfif.rsel1 = SW[9:5];
assign rfif.rsel2 = SW[14:10];
assign rfif.wdat = {29'b0,SW[17:15]};

assign rfif.WEN = ~KEY[3];

assign LEDR[8:5] = rfif.rdat1[3:0];
assign LEDR[13:10] = rfif.rdat2[3:0];
*/

endmodule
